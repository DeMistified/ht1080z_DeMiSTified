
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f0",x"e5",x"c3",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"f0",x"e5",x"c3"),
    14 => (x"48",x"e8",x"d1",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c0",x"eb"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"73",x"1e",x"4f"),
    50 => (x"05",x"a9",x"73",x"81"),
    51 => (x"87",x"f9",x"53",x"72"),
    52 => (x"73",x"1e",x"4f",x"26"),
    53 => (x"02",x"9a",x"72",x"1e"),
    54 => (x"c0",x"87",x"e7",x"c0"),
    55 => (x"72",x"4b",x"c1",x"48"),
    56 => (x"87",x"d1",x"06",x"a9"),
    57 => (x"c9",x"06",x"82",x"72"),
    58 => (x"72",x"83",x"73",x"87"),
    59 => (x"87",x"f4",x"01",x"a9"),
    60 => (x"b2",x"c1",x"87",x"c3"),
    61 => (x"03",x"a9",x"72",x"3a"),
    62 => (x"07",x"80",x"73",x"89"),
    63 => (x"05",x"2b",x"2a",x"c1"),
    64 => (x"4b",x"26",x"87",x"f3"),
    65 => (x"75",x"1e",x"4f",x"26"),
    66 => (x"71",x"4d",x"c4",x"1e"),
    67 => (x"ff",x"04",x"a1",x"b7"),
    68 => (x"c3",x"81",x"c1",x"b9"),
    69 => (x"b7",x"72",x"07",x"bd"),
    70 => (x"ba",x"ff",x"04",x"a2"),
    71 => (x"bd",x"c1",x"82",x"c1"),
    72 => (x"87",x"ee",x"fe",x"07"),
    73 => (x"ff",x"04",x"2d",x"c1"),
    74 => (x"07",x"80",x"c1",x"b8"),
    75 => (x"b9",x"ff",x"04",x"2d"),
    76 => (x"26",x"07",x"81",x"c1"),
    77 => (x"1e",x"4f",x"26",x"4d"),
    78 => (x"66",x"c4",x"4a",x"71"),
    79 => (x"88",x"c1",x"48",x"49"),
    80 => (x"71",x"58",x"a6",x"c8"),
    81 => (x"87",x"d4",x"02",x"99"),
    82 => (x"d4",x"ff",x"48",x"12"),
    83 => (x"66",x"c4",x"78",x"08"),
    84 => (x"88",x"c1",x"48",x"49"),
    85 => (x"71",x"58",x"a6",x"c8"),
    86 => (x"87",x"ec",x"05",x"99"),
    87 => (x"71",x"1e",x"4f",x"26"),
    88 => (x"49",x"66",x"c4",x"4a"),
    89 => (x"c8",x"88",x"c1",x"48"),
    90 => (x"99",x"71",x"58",x"a6"),
    91 => (x"ff",x"87",x"d6",x"02"),
    92 => (x"ff",x"c3",x"48",x"d4"),
    93 => (x"c4",x"52",x"68",x"78"),
    94 => (x"c1",x"48",x"49",x"66"),
    95 => (x"58",x"a6",x"c8",x"88"),
    96 => (x"ea",x"05",x"99",x"71"),
    97 => (x"1e",x"4f",x"26",x"87"),
    98 => (x"d4",x"ff",x"1e",x"73"),
    99 => (x"7b",x"ff",x"c3",x"4b"),
   100 => (x"ff",x"c3",x"4a",x"6b"),
   101 => (x"c8",x"49",x"6b",x"7b"),
   102 => (x"c3",x"b1",x"72",x"32"),
   103 => (x"4a",x"6b",x"7b",x"ff"),
   104 => (x"b2",x"71",x"31",x"c8"),
   105 => (x"6b",x"7b",x"ff",x"c3"),
   106 => (x"72",x"32",x"c8",x"49"),
   107 => (x"c4",x"48",x"71",x"b1"),
   108 => (x"26",x"4d",x"26",x"87"),
   109 => (x"26",x"4b",x"26",x"4c"),
   110 => (x"5b",x"5e",x"0e",x"4f"),
   111 => (x"71",x"0e",x"5d",x"5c"),
   112 => (x"4c",x"d4",x"ff",x"4a"),
   113 => (x"ff",x"c3",x"49",x"72"),
   114 => (x"c3",x"7c",x"71",x"99"),
   115 => (x"05",x"bf",x"e8",x"d1"),
   116 => (x"66",x"d0",x"87",x"c8"),
   117 => (x"d4",x"30",x"c9",x"48"),
   118 => (x"66",x"d0",x"58",x"a6"),
   119 => (x"c3",x"29",x"d8",x"49"),
   120 => (x"7c",x"71",x"99",x"ff"),
   121 => (x"d0",x"49",x"66",x"d0"),
   122 => (x"99",x"ff",x"c3",x"29"),
   123 => (x"66",x"d0",x"7c",x"71"),
   124 => (x"c3",x"29",x"c8",x"49"),
   125 => (x"7c",x"71",x"99",x"ff"),
   126 => (x"c3",x"49",x"66",x"d0"),
   127 => (x"7c",x"71",x"99",x"ff"),
   128 => (x"29",x"d0",x"49",x"72"),
   129 => (x"71",x"99",x"ff",x"c3"),
   130 => (x"c9",x"4b",x"6c",x"7c"),
   131 => (x"c3",x"4d",x"ff",x"f0"),
   132 => (x"d0",x"05",x"ab",x"ff"),
   133 => (x"7c",x"ff",x"c3",x"87"),
   134 => (x"8d",x"c1",x"4b",x"6c"),
   135 => (x"c3",x"87",x"c6",x"02"),
   136 => (x"f0",x"02",x"ab",x"ff"),
   137 => (x"fe",x"48",x"73",x"87"),
   138 => (x"c0",x"1e",x"87",x"c7"),
   139 => (x"48",x"d4",x"ff",x"49"),
   140 => (x"c1",x"78",x"ff",x"c3"),
   141 => (x"b7",x"c8",x"c3",x"81"),
   142 => (x"87",x"f1",x"04",x"a9"),
   143 => (x"73",x"1e",x"4f",x"26"),
   144 => (x"c4",x"87",x"e7",x"1e"),
   145 => (x"c0",x"4b",x"df",x"f8"),
   146 => (x"f0",x"ff",x"c0",x"1e"),
   147 => (x"fd",x"49",x"f7",x"c1"),
   148 => (x"86",x"c4",x"87",x"e7"),
   149 => (x"c0",x"05",x"a8",x"c1"),
   150 => (x"d4",x"ff",x"87",x"ea"),
   151 => (x"78",x"ff",x"c3",x"48"),
   152 => (x"c0",x"c0",x"c0",x"c1"),
   153 => (x"c0",x"1e",x"c0",x"c0"),
   154 => (x"e9",x"c1",x"f0",x"e1"),
   155 => (x"87",x"c9",x"fd",x"49"),
   156 => (x"98",x"70",x"86",x"c4"),
   157 => (x"ff",x"87",x"ca",x"05"),
   158 => (x"ff",x"c3",x"48",x"d4"),
   159 => (x"cb",x"48",x"c1",x"78"),
   160 => (x"87",x"e6",x"fe",x"87"),
   161 => (x"fe",x"05",x"8b",x"c1"),
   162 => (x"48",x"c0",x"87",x"fd"),
   163 => (x"1e",x"87",x"e6",x"fc"),
   164 => (x"d4",x"ff",x"1e",x"73"),
   165 => (x"78",x"ff",x"c3",x"48"),
   166 => (x"1e",x"c0",x"4b",x"d3"),
   167 => (x"c1",x"f0",x"ff",x"c0"),
   168 => (x"d4",x"fc",x"49",x"c1"),
   169 => (x"70",x"86",x"c4",x"87"),
   170 => (x"87",x"ca",x"05",x"98"),
   171 => (x"c3",x"48",x"d4",x"ff"),
   172 => (x"48",x"c1",x"78",x"ff"),
   173 => (x"f1",x"fd",x"87",x"cb"),
   174 => (x"05",x"8b",x"c1",x"87"),
   175 => (x"c0",x"87",x"db",x"ff"),
   176 => (x"87",x"f1",x"fb",x"48"),
   177 => (x"5c",x"5b",x"5e",x"0e"),
   178 => (x"4c",x"d4",x"ff",x"0e"),
   179 => (x"c6",x"87",x"db",x"fd"),
   180 => (x"e1",x"c0",x"1e",x"ea"),
   181 => (x"49",x"c8",x"c1",x"f0"),
   182 => (x"c4",x"87",x"de",x"fb"),
   183 => (x"02",x"a8",x"c1",x"86"),
   184 => (x"ea",x"fe",x"87",x"c8"),
   185 => (x"c1",x"48",x"c0",x"87"),
   186 => (x"da",x"fa",x"87",x"e2"),
   187 => (x"cf",x"49",x"70",x"87"),
   188 => (x"c6",x"99",x"ff",x"ff"),
   189 => (x"c8",x"02",x"a9",x"ea"),
   190 => (x"87",x"d3",x"fe",x"87"),
   191 => (x"cb",x"c1",x"48",x"c0"),
   192 => (x"7c",x"ff",x"c3",x"87"),
   193 => (x"fc",x"4b",x"f1",x"c0"),
   194 => (x"98",x"70",x"87",x"f4"),
   195 => (x"87",x"eb",x"c0",x"02"),
   196 => (x"ff",x"c0",x"1e",x"c0"),
   197 => (x"49",x"fa",x"c1",x"f0"),
   198 => (x"c4",x"87",x"de",x"fa"),
   199 => (x"05",x"98",x"70",x"86"),
   200 => (x"ff",x"c3",x"87",x"d9"),
   201 => (x"c3",x"49",x"6c",x"7c"),
   202 => (x"7c",x"7c",x"7c",x"ff"),
   203 => (x"99",x"c0",x"c1",x"7c"),
   204 => (x"c1",x"87",x"c4",x"02"),
   205 => (x"c0",x"87",x"d5",x"48"),
   206 => (x"c2",x"87",x"d1",x"48"),
   207 => (x"87",x"c4",x"05",x"ab"),
   208 => (x"87",x"c8",x"48",x"c0"),
   209 => (x"fe",x"05",x"8b",x"c1"),
   210 => (x"48",x"c0",x"87",x"fd"),
   211 => (x"1e",x"87",x"e4",x"f9"),
   212 => (x"d1",x"c3",x"1e",x"73"),
   213 => (x"78",x"c1",x"48",x"e8"),
   214 => (x"d0",x"ff",x"4b",x"c7"),
   215 => (x"fb",x"78",x"c2",x"48"),
   216 => (x"d0",x"ff",x"87",x"c8"),
   217 => (x"c0",x"78",x"c3",x"48"),
   218 => (x"d0",x"e5",x"c0",x"1e"),
   219 => (x"f9",x"49",x"c0",x"c1"),
   220 => (x"86",x"c4",x"87",x"c7"),
   221 => (x"c1",x"05",x"a8",x"c1"),
   222 => (x"ab",x"c2",x"4b",x"87"),
   223 => (x"c0",x"87",x"c5",x"05"),
   224 => (x"87",x"f9",x"c0",x"48"),
   225 => (x"ff",x"05",x"8b",x"c1"),
   226 => (x"f7",x"fc",x"87",x"d0"),
   227 => (x"ec",x"d1",x"c3",x"87"),
   228 => (x"05",x"98",x"70",x"58"),
   229 => (x"1e",x"c1",x"87",x"cd"),
   230 => (x"c1",x"f0",x"ff",x"c0"),
   231 => (x"d8",x"f8",x"49",x"d0"),
   232 => (x"ff",x"86",x"c4",x"87"),
   233 => (x"ff",x"c3",x"48",x"d4"),
   234 => (x"87",x"de",x"c4",x"78"),
   235 => (x"58",x"f0",x"d1",x"c3"),
   236 => (x"c2",x"48",x"d0",x"ff"),
   237 => (x"48",x"d4",x"ff",x"78"),
   238 => (x"c1",x"78",x"ff",x"c3"),
   239 => (x"87",x"f5",x"f7",x"48"),
   240 => (x"5c",x"5b",x"5e",x"0e"),
   241 => (x"4a",x"71",x"0e",x"5d"),
   242 => (x"ff",x"4d",x"ff",x"c3"),
   243 => (x"7c",x"75",x"4c",x"d4"),
   244 => (x"c4",x"48",x"d0",x"ff"),
   245 => (x"7c",x"75",x"78",x"c3"),
   246 => (x"ff",x"c0",x"1e",x"72"),
   247 => (x"49",x"d8",x"c1",x"f0"),
   248 => (x"c4",x"87",x"d6",x"f7"),
   249 => (x"02",x"98",x"70",x"86"),
   250 => (x"48",x"c1",x"87",x"c5"),
   251 => (x"75",x"87",x"f0",x"c0"),
   252 => (x"7c",x"fe",x"c3",x"7c"),
   253 => (x"d4",x"1e",x"c0",x"c8"),
   254 => (x"fa",x"f4",x"49",x"66"),
   255 => (x"75",x"86",x"c4",x"87"),
   256 => (x"75",x"7c",x"75",x"7c"),
   257 => (x"e0",x"da",x"d8",x"7c"),
   258 => (x"6c",x"7c",x"75",x"4b"),
   259 => (x"c5",x"05",x"99",x"49"),
   260 => (x"05",x"8b",x"c1",x"87"),
   261 => (x"7c",x"75",x"87",x"f3"),
   262 => (x"c2",x"48",x"d0",x"ff"),
   263 => (x"f6",x"48",x"c0",x"78"),
   264 => (x"5e",x"0e",x"87",x"cf"),
   265 => (x"0e",x"5d",x"5c",x"5b"),
   266 => (x"4c",x"c0",x"4b",x"71"),
   267 => (x"df",x"cd",x"ee",x"c5"),
   268 => (x"48",x"d4",x"ff",x"4a"),
   269 => (x"68",x"78",x"ff",x"c3"),
   270 => (x"a9",x"fe",x"c3",x"49"),
   271 => (x"87",x"fd",x"c0",x"05"),
   272 => (x"9b",x"73",x"4d",x"70"),
   273 => (x"d0",x"87",x"cc",x"02"),
   274 => (x"49",x"73",x"1e",x"66"),
   275 => (x"c4",x"87",x"cf",x"f4"),
   276 => (x"ff",x"87",x"d6",x"86"),
   277 => (x"d1",x"c4",x"48",x"d0"),
   278 => (x"7d",x"ff",x"c3",x"78"),
   279 => (x"c1",x"48",x"66",x"d0"),
   280 => (x"58",x"a6",x"d4",x"88"),
   281 => (x"f0",x"05",x"98",x"70"),
   282 => (x"48",x"d4",x"ff",x"87"),
   283 => (x"78",x"78",x"ff",x"c3"),
   284 => (x"c5",x"05",x"9b",x"73"),
   285 => (x"48",x"d0",x"ff",x"87"),
   286 => (x"4a",x"c1",x"78",x"d0"),
   287 => (x"05",x"8a",x"c1",x"4c"),
   288 => (x"74",x"87",x"ee",x"fe"),
   289 => (x"87",x"e9",x"f4",x"48"),
   290 => (x"71",x"1e",x"73",x"1e"),
   291 => (x"ff",x"4b",x"c0",x"4a"),
   292 => (x"ff",x"c3",x"48",x"d4"),
   293 => (x"48",x"d0",x"ff",x"78"),
   294 => (x"ff",x"78",x"c3",x"c4"),
   295 => (x"ff",x"c3",x"48",x"d4"),
   296 => (x"c0",x"1e",x"72",x"78"),
   297 => (x"d1",x"c1",x"f0",x"ff"),
   298 => (x"87",x"cd",x"f4",x"49"),
   299 => (x"98",x"70",x"86",x"c4"),
   300 => (x"c8",x"87",x"d2",x"05"),
   301 => (x"66",x"cc",x"1e",x"c0"),
   302 => (x"87",x"e6",x"fd",x"49"),
   303 => (x"4b",x"70",x"86",x"c4"),
   304 => (x"c2",x"48",x"d0",x"ff"),
   305 => (x"f3",x"48",x"73",x"78"),
   306 => (x"5e",x"0e",x"87",x"eb"),
   307 => (x"0e",x"5d",x"5c",x"5b"),
   308 => (x"ff",x"c0",x"1e",x"c0"),
   309 => (x"49",x"c9",x"c1",x"f0"),
   310 => (x"d2",x"87",x"de",x"f3"),
   311 => (x"f0",x"d1",x"c3",x"1e"),
   312 => (x"87",x"fe",x"fc",x"49"),
   313 => (x"4c",x"c0",x"86",x"c8"),
   314 => (x"b7",x"d2",x"84",x"c1"),
   315 => (x"87",x"f8",x"04",x"ac"),
   316 => (x"97",x"f0",x"d1",x"c3"),
   317 => (x"c0",x"c3",x"49",x"bf"),
   318 => (x"a9",x"c0",x"c1",x"99"),
   319 => (x"87",x"e7",x"c0",x"05"),
   320 => (x"97",x"f7",x"d1",x"c3"),
   321 => (x"31",x"d0",x"49",x"bf"),
   322 => (x"97",x"f8",x"d1",x"c3"),
   323 => (x"32",x"c8",x"4a",x"bf"),
   324 => (x"d1",x"c3",x"b1",x"72"),
   325 => (x"4a",x"bf",x"97",x"f9"),
   326 => (x"cf",x"4c",x"71",x"b1"),
   327 => (x"9c",x"ff",x"ff",x"ff"),
   328 => (x"34",x"ca",x"84",x"c1"),
   329 => (x"c3",x"87",x"e7",x"c1"),
   330 => (x"bf",x"97",x"f9",x"d1"),
   331 => (x"c6",x"31",x"c1",x"49"),
   332 => (x"fa",x"d1",x"c3",x"99"),
   333 => (x"c7",x"4a",x"bf",x"97"),
   334 => (x"b1",x"72",x"2a",x"b7"),
   335 => (x"97",x"f5",x"d1",x"c3"),
   336 => (x"cf",x"4d",x"4a",x"bf"),
   337 => (x"f6",x"d1",x"c3",x"9d"),
   338 => (x"c3",x"4a",x"bf",x"97"),
   339 => (x"c3",x"32",x"ca",x"9a"),
   340 => (x"bf",x"97",x"f7",x"d1"),
   341 => (x"73",x"33",x"c2",x"4b"),
   342 => (x"f8",x"d1",x"c3",x"b2"),
   343 => (x"c3",x"4b",x"bf",x"97"),
   344 => (x"b7",x"c6",x"9b",x"c0"),
   345 => (x"c2",x"b2",x"73",x"2b"),
   346 => (x"71",x"48",x"c1",x"81"),
   347 => (x"c1",x"49",x"70",x"30"),
   348 => (x"70",x"30",x"75",x"48"),
   349 => (x"c1",x"4c",x"72",x"4d"),
   350 => (x"c8",x"94",x"71",x"84"),
   351 => (x"06",x"ad",x"b7",x"c0"),
   352 => (x"34",x"c1",x"87",x"cc"),
   353 => (x"c0",x"c8",x"2d",x"b7"),
   354 => (x"ff",x"01",x"ad",x"b7"),
   355 => (x"48",x"74",x"87",x"f4"),
   356 => (x"0e",x"87",x"de",x"f0"),
   357 => (x"5d",x"5c",x"5b",x"5e"),
   358 => (x"c3",x"86",x"f8",x"0e"),
   359 => (x"c0",x"48",x"d6",x"da"),
   360 => (x"ce",x"d2",x"c3",x"78"),
   361 => (x"fb",x"49",x"c0",x"1e"),
   362 => (x"86",x"c4",x"87",x"de"),
   363 => (x"c5",x"05",x"98",x"70"),
   364 => (x"c9",x"48",x"c0",x"87"),
   365 => (x"4d",x"c0",x"87",x"ce"),
   366 => (x"fa",x"c0",x"7e",x"c1"),
   367 => (x"c3",x"49",x"bf",x"e1"),
   368 => (x"71",x"4a",x"c4",x"d3"),
   369 => (x"e1",x"ea",x"4b",x"c8"),
   370 => (x"05",x"98",x"70",x"87"),
   371 => (x"7e",x"c0",x"87",x"c2"),
   372 => (x"bf",x"dd",x"fa",x"c0"),
   373 => (x"e0",x"d3",x"c3",x"49"),
   374 => (x"4b",x"c8",x"71",x"4a"),
   375 => (x"70",x"87",x"cb",x"ea"),
   376 => (x"87",x"c2",x"05",x"98"),
   377 => (x"02",x"6e",x"7e",x"c0"),
   378 => (x"c3",x"87",x"fd",x"c0"),
   379 => (x"4d",x"bf",x"d4",x"d9"),
   380 => (x"9f",x"cc",x"da",x"c3"),
   381 => (x"c5",x"48",x"7e",x"bf"),
   382 => (x"05",x"a8",x"ea",x"d6"),
   383 => (x"d9",x"c3",x"87",x"c7"),
   384 => (x"ce",x"4d",x"bf",x"d4"),
   385 => (x"ca",x"48",x"6e",x"87"),
   386 => (x"02",x"a8",x"d5",x"e9"),
   387 => (x"48",x"c0",x"87",x"c5"),
   388 => (x"c3",x"87",x"f1",x"c7"),
   389 => (x"75",x"1e",x"ce",x"d2"),
   390 => (x"87",x"ec",x"f9",x"49"),
   391 => (x"98",x"70",x"86",x"c4"),
   392 => (x"c0",x"87",x"c5",x"05"),
   393 => (x"87",x"dc",x"c7",x"48"),
   394 => (x"bf",x"dd",x"fa",x"c0"),
   395 => (x"e0",x"d3",x"c3",x"49"),
   396 => (x"4b",x"c8",x"71",x"4a"),
   397 => (x"70",x"87",x"f3",x"e8"),
   398 => (x"87",x"c8",x"05",x"98"),
   399 => (x"48",x"d6",x"da",x"c3"),
   400 => (x"87",x"da",x"78",x"c1"),
   401 => (x"bf",x"e1",x"fa",x"c0"),
   402 => (x"c4",x"d3",x"c3",x"49"),
   403 => (x"4b",x"c8",x"71",x"4a"),
   404 => (x"70",x"87",x"d7",x"e8"),
   405 => (x"c5",x"c0",x"02",x"98"),
   406 => (x"c6",x"48",x"c0",x"87"),
   407 => (x"da",x"c3",x"87",x"e6"),
   408 => (x"49",x"bf",x"97",x"cc"),
   409 => (x"05",x"a9",x"d5",x"c1"),
   410 => (x"c3",x"87",x"cd",x"c0"),
   411 => (x"bf",x"97",x"cd",x"da"),
   412 => (x"a9",x"ea",x"c2",x"49"),
   413 => (x"87",x"c5",x"c0",x"02"),
   414 => (x"c7",x"c6",x"48",x"c0"),
   415 => (x"ce",x"d2",x"c3",x"87"),
   416 => (x"48",x"7e",x"bf",x"97"),
   417 => (x"02",x"a8",x"e9",x"c3"),
   418 => (x"6e",x"87",x"ce",x"c0"),
   419 => (x"a8",x"eb",x"c3",x"48"),
   420 => (x"87",x"c5",x"c0",x"02"),
   421 => (x"eb",x"c5",x"48",x"c0"),
   422 => (x"d9",x"d2",x"c3",x"87"),
   423 => (x"99",x"49",x"bf",x"97"),
   424 => (x"87",x"cc",x"c0",x"05"),
   425 => (x"97",x"da",x"d2",x"c3"),
   426 => (x"a9",x"c2",x"49",x"bf"),
   427 => (x"87",x"c5",x"c0",x"02"),
   428 => (x"cf",x"c5",x"48",x"c0"),
   429 => (x"db",x"d2",x"c3",x"87"),
   430 => (x"c3",x"48",x"bf",x"97"),
   431 => (x"70",x"58",x"d2",x"da"),
   432 => (x"88",x"c1",x"48",x"4c"),
   433 => (x"58",x"d6",x"da",x"c3"),
   434 => (x"97",x"dc",x"d2",x"c3"),
   435 => (x"81",x"75",x"49",x"bf"),
   436 => (x"97",x"dd",x"d2",x"c3"),
   437 => (x"32",x"c8",x"4a",x"bf"),
   438 => (x"c3",x"7e",x"a1",x"72"),
   439 => (x"6e",x"48",x"e3",x"de"),
   440 => (x"de",x"d2",x"c3",x"78"),
   441 => (x"c8",x"48",x"bf",x"97"),
   442 => (x"da",x"c3",x"58",x"a6"),
   443 => (x"c2",x"02",x"bf",x"d6"),
   444 => (x"fa",x"c0",x"87",x"d4"),
   445 => (x"c3",x"49",x"bf",x"dd"),
   446 => (x"71",x"4a",x"e0",x"d3"),
   447 => (x"e9",x"e5",x"4b",x"c8"),
   448 => (x"02",x"98",x"70",x"87"),
   449 => (x"c0",x"87",x"c5",x"c0"),
   450 => (x"87",x"f8",x"c3",x"48"),
   451 => (x"bf",x"ce",x"da",x"c3"),
   452 => (x"f7",x"de",x"c3",x"4c"),
   453 => (x"f3",x"d2",x"c3",x"5c"),
   454 => (x"c8",x"49",x"bf",x"97"),
   455 => (x"f2",x"d2",x"c3",x"31"),
   456 => (x"a1",x"4a",x"bf",x"97"),
   457 => (x"f4",x"d2",x"c3",x"49"),
   458 => (x"d0",x"4a",x"bf",x"97"),
   459 => (x"49",x"a1",x"72",x"32"),
   460 => (x"97",x"f5",x"d2",x"c3"),
   461 => (x"32",x"d8",x"4a",x"bf"),
   462 => (x"c4",x"49",x"a1",x"72"),
   463 => (x"de",x"c3",x"91",x"66"),
   464 => (x"c3",x"81",x"bf",x"e3"),
   465 => (x"c3",x"59",x"eb",x"de"),
   466 => (x"bf",x"97",x"fb",x"d2"),
   467 => (x"c3",x"32",x"c8",x"4a"),
   468 => (x"bf",x"97",x"fa",x"d2"),
   469 => (x"c3",x"4a",x"a2",x"4b"),
   470 => (x"bf",x"97",x"fc",x"d2"),
   471 => (x"73",x"33",x"d0",x"4b"),
   472 => (x"d2",x"c3",x"4a",x"a2"),
   473 => (x"4b",x"bf",x"97",x"fd"),
   474 => (x"33",x"d8",x"9b",x"cf"),
   475 => (x"c3",x"4a",x"a2",x"73"),
   476 => (x"c3",x"5a",x"ef",x"de"),
   477 => (x"4a",x"bf",x"eb",x"de"),
   478 => (x"92",x"74",x"8a",x"c2"),
   479 => (x"48",x"ef",x"de",x"c3"),
   480 => (x"c1",x"78",x"a1",x"72"),
   481 => (x"d2",x"c3",x"87",x"ca"),
   482 => (x"49",x"bf",x"97",x"e0"),
   483 => (x"d2",x"c3",x"31",x"c8"),
   484 => (x"4a",x"bf",x"97",x"df"),
   485 => (x"da",x"c3",x"49",x"a1"),
   486 => (x"da",x"c3",x"59",x"de"),
   487 => (x"c5",x"49",x"bf",x"da"),
   488 => (x"81",x"ff",x"c7",x"31"),
   489 => (x"de",x"c3",x"29",x"c9"),
   490 => (x"d2",x"c3",x"59",x"f7"),
   491 => (x"4a",x"bf",x"97",x"e5"),
   492 => (x"d2",x"c3",x"32",x"c8"),
   493 => (x"4b",x"bf",x"97",x"e4"),
   494 => (x"66",x"c4",x"4a",x"a2"),
   495 => (x"c3",x"82",x"6e",x"92"),
   496 => (x"c3",x"5a",x"f3",x"de"),
   497 => (x"c0",x"48",x"eb",x"de"),
   498 => (x"e7",x"de",x"c3",x"78"),
   499 => (x"78",x"a1",x"72",x"48"),
   500 => (x"48",x"f7",x"de",x"c3"),
   501 => (x"bf",x"eb",x"de",x"c3"),
   502 => (x"fb",x"de",x"c3",x"78"),
   503 => (x"ef",x"de",x"c3",x"48"),
   504 => (x"da",x"c3",x"78",x"bf"),
   505 => (x"c0",x"02",x"bf",x"d6"),
   506 => (x"48",x"74",x"87",x"c9"),
   507 => (x"7e",x"70",x"30",x"c4"),
   508 => (x"c3",x"87",x"c9",x"c0"),
   509 => (x"48",x"bf",x"f3",x"de"),
   510 => (x"7e",x"70",x"30",x"c4"),
   511 => (x"48",x"da",x"da",x"c3"),
   512 => (x"48",x"c1",x"78",x"6e"),
   513 => (x"4d",x"26",x"8e",x"f8"),
   514 => (x"4b",x"26",x"4c",x"26"),
   515 => (x"5e",x"0e",x"4f",x"26"),
   516 => (x"0e",x"5d",x"5c",x"5b"),
   517 => (x"da",x"c3",x"4a",x"71"),
   518 => (x"cb",x"02",x"bf",x"d6"),
   519 => (x"c7",x"4b",x"72",x"87"),
   520 => (x"c1",x"4c",x"72",x"2b"),
   521 => (x"87",x"c9",x"9c",x"ff"),
   522 => (x"2b",x"c8",x"4b",x"72"),
   523 => (x"ff",x"c3",x"4c",x"72"),
   524 => (x"e3",x"de",x"c3",x"9c"),
   525 => (x"fa",x"c0",x"83",x"bf"),
   526 => (x"02",x"ab",x"bf",x"d9"),
   527 => (x"fa",x"c0",x"87",x"d9"),
   528 => (x"d2",x"c3",x"5b",x"dd"),
   529 => (x"49",x"73",x"1e",x"ce"),
   530 => (x"c4",x"87",x"fd",x"f0"),
   531 => (x"05",x"98",x"70",x"86"),
   532 => (x"48",x"c0",x"87",x"c5"),
   533 => (x"c3",x"87",x"e6",x"c0"),
   534 => (x"02",x"bf",x"d6",x"da"),
   535 => (x"49",x"74",x"87",x"d2"),
   536 => (x"d2",x"c3",x"91",x"c4"),
   537 => (x"4d",x"69",x"81",x"ce"),
   538 => (x"ff",x"ff",x"ff",x"cf"),
   539 => (x"87",x"cb",x"9d",x"ff"),
   540 => (x"91",x"c2",x"49",x"74"),
   541 => (x"81",x"ce",x"d2",x"c3"),
   542 => (x"75",x"4d",x"69",x"9f"),
   543 => (x"87",x"c6",x"fe",x"48"),
   544 => (x"5c",x"5b",x"5e",x"0e"),
   545 => (x"71",x"1e",x"0e",x"5d"),
   546 => (x"c1",x"1e",x"c0",x"4d"),
   547 => (x"87",x"ed",x"d0",x"49"),
   548 => (x"4c",x"70",x"86",x"c4"),
   549 => (x"c2",x"c1",x"02",x"9c"),
   550 => (x"de",x"da",x"c3",x"87"),
   551 => (x"ff",x"49",x"75",x"4a"),
   552 => (x"70",x"87",x"ec",x"de"),
   553 => (x"f2",x"c0",x"02",x"98"),
   554 => (x"75",x"4a",x"74",x"87"),
   555 => (x"ff",x"4b",x"cb",x"49"),
   556 => (x"70",x"87",x"d1",x"df"),
   557 => (x"e2",x"c0",x"02",x"98"),
   558 => (x"74",x"1e",x"c0",x"87"),
   559 => (x"87",x"c7",x"02",x"9c"),
   560 => (x"c0",x"48",x"a6",x"c4"),
   561 => (x"c4",x"87",x"c5",x"78"),
   562 => (x"78",x"c1",x"48",x"a6"),
   563 => (x"cf",x"49",x"66",x"c4"),
   564 => (x"86",x"c4",x"87",x"eb"),
   565 => (x"05",x"9c",x"4c",x"70"),
   566 => (x"74",x"87",x"fe",x"fe"),
   567 => (x"e5",x"fc",x"26",x"48"),
   568 => (x"5b",x"5e",x"0e",x"87"),
   569 => (x"1e",x"0e",x"5d",x"5c"),
   570 => (x"05",x"9b",x"4b",x"71"),
   571 => (x"48",x"c0",x"87",x"c5"),
   572 => (x"c8",x"87",x"e5",x"c1"),
   573 => (x"7d",x"c0",x"4d",x"a3"),
   574 => (x"c7",x"02",x"66",x"d4"),
   575 => (x"97",x"66",x"d4",x"87"),
   576 => (x"87",x"c5",x"05",x"bf"),
   577 => (x"cf",x"c1",x"48",x"c0"),
   578 => (x"49",x"66",x"d4",x"87"),
   579 => (x"70",x"87",x"f1",x"fd"),
   580 => (x"c1",x"02",x"9c",x"4c"),
   581 => (x"a4",x"dc",x"87",x"c0"),
   582 => (x"da",x"7d",x"69",x"49"),
   583 => (x"a3",x"c4",x"49",x"a4"),
   584 => (x"7a",x"69",x"9f",x"4a"),
   585 => (x"bf",x"d6",x"da",x"c3"),
   586 => (x"d4",x"87",x"d2",x"02"),
   587 => (x"69",x"9f",x"49",x"a4"),
   588 => (x"ff",x"ff",x"c0",x"49"),
   589 => (x"d0",x"48",x"71",x"99"),
   590 => (x"c2",x"7e",x"70",x"30"),
   591 => (x"6e",x"7e",x"c0",x"87"),
   592 => (x"80",x"6a",x"48",x"49"),
   593 => (x"7b",x"c0",x"7a",x"70"),
   594 => (x"6a",x"49",x"a3",x"cc"),
   595 => (x"49",x"a3",x"d0",x"79"),
   596 => (x"48",x"c1",x"79",x"c0"),
   597 => (x"48",x"c0",x"87",x"c2"),
   598 => (x"87",x"ea",x"fa",x"26"),
   599 => (x"5c",x"5b",x"5e",x"0e"),
   600 => (x"4c",x"71",x"0e",x"5d"),
   601 => (x"ca",x"c1",x"02",x"9c"),
   602 => (x"49",x"a4",x"c8",x"87"),
   603 => (x"c2",x"c1",x"02",x"69"),
   604 => (x"4a",x"66",x"d0",x"87"),
   605 => (x"d4",x"82",x"49",x"6c"),
   606 => (x"66",x"d0",x"5a",x"a6"),
   607 => (x"da",x"c3",x"b9",x"4d"),
   608 => (x"ff",x"4a",x"bf",x"d2"),
   609 => (x"71",x"99",x"72",x"ba"),
   610 => (x"e4",x"c0",x"02",x"99"),
   611 => (x"4b",x"a4",x"c4",x"87"),
   612 => (x"f9",x"f9",x"49",x"6b"),
   613 => (x"c3",x"7b",x"70",x"87"),
   614 => (x"49",x"bf",x"ce",x"da"),
   615 => (x"7c",x"71",x"81",x"6c"),
   616 => (x"da",x"c3",x"b9",x"75"),
   617 => (x"ff",x"4a",x"bf",x"d2"),
   618 => (x"71",x"99",x"72",x"ba"),
   619 => (x"dc",x"ff",x"05",x"99"),
   620 => (x"f9",x"7c",x"75",x"87"),
   621 => (x"73",x"1e",x"87",x"d0"),
   622 => (x"9b",x"4b",x"71",x"1e"),
   623 => (x"c8",x"87",x"c7",x"02"),
   624 => (x"05",x"69",x"49",x"a3"),
   625 => (x"48",x"c0",x"87",x"c5"),
   626 => (x"c3",x"87",x"f7",x"c0"),
   627 => (x"4a",x"bf",x"e7",x"de"),
   628 => (x"69",x"49",x"a3",x"c4"),
   629 => (x"c3",x"89",x"c2",x"49"),
   630 => (x"91",x"bf",x"ce",x"da"),
   631 => (x"c3",x"4a",x"a2",x"71"),
   632 => (x"49",x"bf",x"d2",x"da"),
   633 => (x"a2",x"71",x"99",x"6b"),
   634 => (x"dd",x"fa",x"c0",x"4a"),
   635 => (x"1e",x"66",x"c8",x"5a"),
   636 => (x"d3",x"ea",x"49",x"72"),
   637 => (x"70",x"86",x"c4",x"87"),
   638 => (x"87",x"c4",x"05",x"98"),
   639 => (x"87",x"c2",x"48",x"c0"),
   640 => (x"c5",x"f8",x"48",x"c1"),
   641 => (x"1e",x"73",x"1e",x"87"),
   642 => (x"02",x"9b",x"4b",x"71"),
   643 => (x"a3",x"c8",x"87",x"c7"),
   644 => (x"c5",x"05",x"69",x"49"),
   645 => (x"c0",x"48",x"c0",x"87"),
   646 => (x"de",x"c3",x"87",x"f7"),
   647 => (x"c4",x"4a",x"bf",x"e7"),
   648 => (x"49",x"69",x"49",x"a3"),
   649 => (x"da",x"c3",x"89",x"c2"),
   650 => (x"71",x"91",x"bf",x"ce"),
   651 => (x"da",x"c3",x"4a",x"a2"),
   652 => (x"6b",x"49",x"bf",x"d2"),
   653 => (x"4a",x"a2",x"71",x"99"),
   654 => (x"5a",x"dd",x"fa",x"c0"),
   655 => (x"72",x"1e",x"66",x"c8"),
   656 => (x"87",x"fc",x"e5",x"49"),
   657 => (x"98",x"70",x"86",x"c4"),
   658 => (x"c0",x"87",x"c4",x"05"),
   659 => (x"c1",x"87",x"c2",x"48"),
   660 => (x"87",x"f6",x"f6",x"48"),
   661 => (x"5c",x"5b",x"5e",x"0e"),
   662 => (x"71",x"1e",x"0e",x"5d"),
   663 => (x"4c",x"66",x"d4",x"4b"),
   664 => (x"9b",x"73",x"2c",x"c9"),
   665 => (x"87",x"cf",x"c1",x"02"),
   666 => (x"69",x"49",x"a3",x"c8"),
   667 => (x"87",x"c7",x"c1",x"02"),
   668 => (x"d4",x"4d",x"a3",x"d0"),
   669 => (x"da",x"c3",x"7d",x"66"),
   670 => (x"ff",x"49",x"bf",x"d2"),
   671 => (x"99",x"4a",x"6b",x"b9"),
   672 => (x"03",x"ac",x"71",x"7e"),
   673 => (x"7b",x"c0",x"87",x"cd"),
   674 => (x"4a",x"a3",x"cc",x"7d"),
   675 => (x"6a",x"49",x"a3",x"c4"),
   676 => (x"72",x"87",x"c2",x"79"),
   677 => (x"02",x"9c",x"74",x"8c"),
   678 => (x"1e",x"49",x"87",x"dd"),
   679 => (x"fb",x"fa",x"49",x"73"),
   680 => (x"d4",x"86",x"c4",x"87"),
   681 => (x"ff",x"c7",x"49",x"66"),
   682 => (x"87",x"cb",x"02",x"99"),
   683 => (x"1e",x"ce",x"d2",x"c3"),
   684 => (x"c1",x"fc",x"49",x"73"),
   685 => (x"26",x"86",x"c4",x"87"),
   686 => (x"0e",x"87",x"cb",x"f5"),
   687 => (x"5d",x"5c",x"5b",x"5e"),
   688 => (x"d0",x"86",x"f0",x"0e"),
   689 => (x"e4",x"c0",x"59",x"a6"),
   690 => (x"66",x"cc",x"4b",x"66"),
   691 => (x"48",x"87",x"ca",x"02"),
   692 => (x"7e",x"70",x"80",x"c8"),
   693 => (x"c5",x"05",x"bf",x"6e"),
   694 => (x"c3",x"48",x"c0",x"87"),
   695 => (x"66",x"cc",x"87",x"ec"),
   696 => (x"73",x"84",x"d0",x"4c"),
   697 => (x"48",x"a6",x"c4",x"49"),
   698 => (x"66",x"c4",x"78",x"6c"),
   699 => (x"6e",x"80",x"c4",x"81"),
   700 => (x"66",x"c8",x"78",x"bf"),
   701 => (x"87",x"c6",x"06",x"a9"),
   702 => (x"89",x"66",x"c4",x"49"),
   703 => (x"b7",x"c0",x"4b",x"71"),
   704 => (x"87",x"c4",x"01",x"ab"),
   705 => (x"87",x"c2",x"c3",x"48"),
   706 => (x"c7",x"48",x"66",x"c4"),
   707 => (x"7e",x"70",x"98",x"ff"),
   708 => (x"c9",x"c1",x"02",x"6e"),
   709 => (x"49",x"c0",x"c8",x"87"),
   710 => (x"4a",x"71",x"89",x"6e"),
   711 => (x"4d",x"ce",x"d2",x"c3"),
   712 => (x"b7",x"73",x"85",x"6e"),
   713 => (x"87",x"c1",x"06",x"aa"),
   714 => (x"48",x"49",x"72",x"4a"),
   715 => (x"70",x"80",x"66",x"c4"),
   716 => (x"49",x"8b",x"72",x"7c"),
   717 => (x"99",x"71",x"8a",x"c1"),
   718 => (x"c0",x"87",x"d9",x"02"),
   719 => (x"15",x"48",x"66",x"e0"),
   720 => (x"66",x"e0",x"c0",x"50"),
   721 => (x"c0",x"80",x"c1",x"48"),
   722 => (x"72",x"58",x"a6",x"e4"),
   723 => (x"71",x"8a",x"c1",x"49"),
   724 => (x"87",x"e7",x"05",x"99"),
   725 => (x"66",x"d0",x"1e",x"c1"),
   726 => (x"87",x"c0",x"f8",x"49"),
   727 => (x"b7",x"c0",x"86",x"c4"),
   728 => (x"e3",x"c1",x"06",x"ab"),
   729 => (x"66",x"e0",x"c0",x"87"),
   730 => (x"b7",x"ff",x"c7",x"4d"),
   731 => (x"e2",x"c0",x"06",x"ab"),
   732 => (x"d0",x"1e",x"75",x"87"),
   733 => (x"fd",x"f8",x"49",x"66"),
   734 => (x"85",x"c0",x"c8",x"87"),
   735 => (x"c0",x"c8",x"48",x"6c"),
   736 => (x"c8",x"7c",x"70",x"80"),
   737 => (x"1e",x"c1",x"8b",x"c0"),
   738 => (x"f7",x"49",x"66",x"d4"),
   739 => (x"86",x"c8",x"87",x"ce"),
   740 => (x"c3",x"87",x"ee",x"c0"),
   741 => (x"d0",x"1e",x"ce",x"d2"),
   742 => (x"d9",x"f8",x"49",x"66"),
   743 => (x"c3",x"86",x"c4",x"87"),
   744 => (x"73",x"4a",x"ce",x"d2"),
   745 => (x"80",x"6c",x"48",x"49"),
   746 => (x"49",x"73",x"7c",x"70"),
   747 => (x"99",x"71",x"8b",x"c1"),
   748 => (x"12",x"87",x"ce",x"02"),
   749 => (x"85",x"c1",x"7d",x"97"),
   750 => (x"8b",x"c1",x"49",x"73"),
   751 => (x"f2",x"05",x"99",x"71"),
   752 => (x"ab",x"b7",x"c0",x"87"),
   753 => (x"87",x"e1",x"fe",x"01"),
   754 => (x"8e",x"f0",x"48",x"c1"),
   755 => (x"0e",x"87",x"f7",x"f0"),
   756 => (x"5d",x"5c",x"5b",x"5e"),
   757 => (x"9b",x"4b",x"71",x"0e"),
   758 => (x"c8",x"87",x"c7",x"02"),
   759 => (x"05",x"6d",x"4d",x"a3"),
   760 => (x"48",x"ff",x"87",x"c5"),
   761 => (x"d0",x"87",x"fd",x"c0"),
   762 => (x"49",x"6c",x"4c",x"a3"),
   763 => (x"05",x"99",x"ff",x"c7"),
   764 => (x"02",x"6c",x"87",x"d8"),
   765 => (x"1e",x"c1",x"87",x"c9"),
   766 => (x"df",x"f5",x"49",x"73"),
   767 => (x"c3",x"86",x"c4",x"87"),
   768 => (x"73",x"1e",x"ce",x"d2"),
   769 => (x"87",x"ee",x"f6",x"49"),
   770 => (x"4a",x"6c",x"86",x"c4"),
   771 => (x"c4",x"04",x"aa",x"6d"),
   772 => (x"cf",x"48",x"ff",x"87"),
   773 => (x"7c",x"a2",x"c1",x"87"),
   774 => (x"ff",x"c7",x"49",x"72"),
   775 => (x"ce",x"d2",x"c3",x"99"),
   776 => (x"48",x"69",x"97",x"81"),
   777 => (x"1e",x"87",x"df",x"ef"),
   778 => (x"4b",x"71",x"1e",x"73"),
   779 => (x"e4",x"c0",x"02",x"9b"),
   780 => (x"fb",x"de",x"c3",x"87"),
   781 => (x"c2",x"4a",x"73",x"5b"),
   782 => (x"ce",x"da",x"c3",x"8a"),
   783 => (x"c3",x"92",x"49",x"bf"),
   784 => (x"48",x"bf",x"e7",x"de"),
   785 => (x"de",x"c3",x"80",x"72"),
   786 => (x"48",x"71",x"58",x"ff"),
   787 => (x"da",x"c3",x"30",x"c4"),
   788 => (x"ed",x"c0",x"58",x"de"),
   789 => (x"f7",x"de",x"c3",x"87"),
   790 => (x"eb",x"de",x"c3",x"48"),
   791 => (x"de",x"c3",x"78",x"bf"),
   792 => (x"de",x"c3",x"48",x"fb"),
   793 => (x"c3",x"78",x"bf",x"ef"),
   794 => (x"02",x"bf",x"d6",x"da"),
   795 => (x"da",x"c3",x"87",x"c9"),
   796 => (x"c4",x"49",x"bf",x"ce"),
   797 => (x"c3",x"87",x"c7",x"31"),
   798 => (x"49",x"bf",x"f3",x"de"),
   799 => (x"da",x"c3",x"31",x"c4"),
   800 => (x"c5",x"ee",x"59",x"de"),
   801 => (x"5b",x"5e",x"0e",x"87"),
   802 => (x"4a",x"71",x"0e",x"5c"),
   803 => (x"9a",x"72",x"4b",x"c0"),
   804 => (x"87",x"e1",x"c0",x"02"),
   805 => (x"9f",x"49",x"a2",x"da"),
   806 => (x"da",x"c3",x"4b",x"69"),
   807 => (x"cf",x"02",x"bf",x"d6"),
   808 => (x"49",x"a2",x"d4",x"87"),
   809 => (x"4c",x"49",x"69",x"9f"),
   810 => (x"9c",x"ff",x"ff",x"c0"),
   811 => (x"87",x"c2",x"34",x"d0"),
   812 => (x"49",x"74",x"4c",x"c0"),
   813 => (x"fd",x"49",x"73",x"b3"),
   814 => (x"cb",x"ed",x"87",x"ed"),
   815 => (x"5b",x"5e",x"0e",x"87"),
   816 => (x"f4",x"0e",x"5d",x"5c"),
   817 => (x"c0",x"4a",x"71",x"86"),
   818 => (x"02",x"9a",x"72",x"7e"),
   819 => (x"d2",x"c3",x"87",x"d8"),
   820 => (x"78",x"c0",x"48",x"ca"),
   821 => (x"48",x"c2",x"d2",x"c3"),
   822 => (x"bf",x"fb",x"de",x"c3"),
   823 => (x"c6",x"d2",x"c3",x"78"),
   824 => (x"f7",x"de",x"c3",x"48"),
   825 => (x"da",x"c3",x"78",x"bf"),
   826 => (x"50",x"c0",x"48",x"eb"),
   827 => (x"bf",x"da",x"da",x"c3"),
   828 => (x"ca",x"d2",x"c3",x"49"),
   829 => (x"aa",x"71",x"4a",x"bf"),
   830 => (x"87",x"ca",x"c4",x"03"),
   831 => (x"99",x"cf",x"49",x"72"),
   832 => (x"87",x"ea",x"c0",x"05"),
   833 => (x"48",x"d9",x"fa",x"c0"),
   834 => (x"bf",x"c2",x"d2",x"c3"),
   835 => (x"ce",x"d2",x"c3",x"78"),
   836 => (x"c2",x"d2",x"c3",x"1e"),
   837 => (x"d2",x"c3",x"49",x"bf"),
   838 => (x"a1",x"c1",x"48",x"c2"),
   839 => (x"dd",x"ff",x"71",x"78"),
   840 => (x"86",x"c4",x"87",x"e6"),
   841 => (x"48",x"d5",x"fa",x"c0"),
   842 => (x"78",x"ce",x"d2",x"c3"),
   843 => (x"fa",x"c0",x"87",x"cc"),
   844 => (x"c0",x"48",x"bf",x"d5"),
   845 => (x"fa",x"c0",x"80",x"e0"),
   846 => (x"d2",x"c3",x"58",x"d9"),
   847 => (x"c1",x"48",x"bf",x"ca"),
   848 => (x"ce",x"d2",x"c3",x"80"),
   849 => (x"0e",x"95",x"27",x"58"),
   850 => (x"97",x"bf",x"00",x"00"),
   851 => (x"02",x"9d",x"4d",x"bf"),
   852 => (x"c3",x"87",x"e3",x"c2"),
   853 => (x"c2",x"02",x"ad",x"e5"),
   854 => (x"fa",x"c0",x"87",x"dc"),
   855 => (x"cb",x"4b",x"bf",x"d5"),
   856 => (x"4c",x"11",x"49",x"a3"),
   857 => (x"c1",x"05",x"ac",x"cf"),
   858 => (x"49",x"75",x"87",x"d2"),
   859 => (x"89",x"c1",x"99",x"df"),
   860 => (x"da",x"c3",x"91",x"cd"),
   861 => (x"a3",x"c1",x"81",x"de"),
   862 => (x"c3",x"51",x"12",x"4a"),
   863 => (x"51",x"12",x"4a",x"a3"),
   864 => (x"12",x"4a",x"a3",x"c5"),
   865 => (x"4a",x"a3",x"c7",x"51"),
   866 => (x"a3",x"c9",x"51",x"12"),
   867 => (x"ce",x"51",x"12",x"4a"),
   868 => (x"51",x"12",x"4a",x"a3"),
   869 => (x"12",x"4a",x"a3",x"d0"),
   870 => (x"4a",x"a3",x"d2",x"51"),
   871 => (x"a3",x"d4",x"51",x"12"),
   872 => (x"d6",x"51",x"12",x"4a"),
   873 => (x"51",x"12",x"4a",x"a3"),
   874 => (x"12",x"4a",x"a3",x"d8"),
   875 => (x"4a",x"a3",x"dc",x"51"),
   876 => (x"a3",x"de",x"51",x"12"),
   877 => (x"c1",x"51",x"12",x"4a"),
   878 => (x"87",x"fa",x"c0",x"7e"),
   879 => (x"99",x"c8",x"49",x"74"),
   880 => (x"87",x"eb",x"c0",x"05"),
   881 => (x"99",x"d0",x"49",x"74"),
   882 => (x"dc",x"87",x"d1",x"05"),
   883 => (x"cb",x"c0",x"02",x"66"),
   884 => (x"dc",x"49",x"73",x"87"),
   885 => (x"98",x"70",x"0f",x"66"),
   886 => (x"87",x"d3",x"c0",x"02"),
   887 => (x"c6",x"c0",x"05",x"6e"),
   888 => (x"de",x"da",x"c3",x"87"),
   889 => (x"c0",x"50",x"c0",x"48"),
   890 => (x"48",x"bf",x"d5",x"fa"),
   891 => (x"c3",x"87",x"e1",x"c2"),
   892 => (x"c0",x"48",x"eb",x"da"),
   893 => (x"da",x"c3",x"7e",x"50"),
   894 => (x"c3",x"49",x"bf",x"da"),
   895 => (x"4a",x"bf",x"ca",x"d2"),
   896 => (x"fb",x"04",x"aa",x"71"),
   897 => (x"de",x"c3",x"87",x"f6"),
   898 => (x"c0",x"05",x"bf",x"fb"),
   899 => (x"da",x"c3",x"87",x"c8"),
   900 => (x"c1",x"02",x"bf",x"d6"),
   901 => (x"d2",x"c3",x"87",x"f8"),
   902 => (x"e7",x"49",x"bf",x"c6"),
   903 => (x"49",x"70",x"87",x"f0"),
   904 => (x"59",x"ca",x"d2",x"c3"),
   905 => (x"c3",x"48",x"a6",x"c4"),
   906 => (x"78",x"bf",x"c6",x"d2"),
   907 => (x"bf",x"d6",x"da",x"c3"),
   908 => (x"87",x"d8",x"c0",x"02"),
   909 => (x"cf",x"49",x"66",x"c4"),
   910 => (x"f8",x"ff",x"ff",x"ff"),
   911 => (x"c0",x"02",x"a9",x"99"),
   912 => (x"4c",x"c0",x"87",x"c5"),
   913 => (x"c1",x"87",x"e1",x"c0"),
   914 => (x"87",x"dc",x"c0",x"4c"),
   915 => (x"cf",x"49",x"66",x"c4"),
   916 => (x"a9",x"99",x"f8",x"ff"),
   917 => (x"87",x"c8",x"c0",x"02"),
   918 => (x"c0",x"48",x"a6",x"c8"),
   919 => (x"87",x"c5",x"c0",x"78"),
   920 => (x"c1",x"48",x"a6",x"c8"),
   921 => (x"4c",x"66",x"c8",x"78"),
   922 => (x"c0",x"05",x"9c",x"74"),
   923 => (x"66",x"c4",x"87",x"e0"),
   924 => (x"c3",x"89",x"c2",x"49"),
   925 => (x"4a",x"bf",x"ce",x"da"),
   926 => (x"e7",x"de",x"c3",x"91"),
   927 => (x"d2",x"c3",x"4a",x"bf"),
   928 => (x"a1",x"72",x"48",x"c2"),
   929 => (x"ca",x"d2",x"c3",x"78"),
   930 => (x"f9",x"78",x"c0",x"48"),
   931 => (x"48",x"c0",x"87",x"de"),
   932 => (x"f1",x"e5",x"8e",x"f4"),
   933 => (x"00",x"00",x"00",x"87"),
   934 => (x"ff",x"ff",x"ff",x"00"),
   935 => (x"00",x"0e",x"a5",x"ff"),
   936 => (x"00",x"0e",x"ae",x"00"),
   937 => (x"54",x"41",x"46",x"00"),
   938 => (x"20",x"20",x"32",x"33"),
   939 => (x"41",x"46",x"00",x"20"),
   940 => (x"20",x"36",x"31",x"54"),
   941 => (x"1e",x"00",x"20",x"20"),
   942 => (x"bf",x"c0",x"df",x"c3"),
   943 => (x"05",x"a8",x"dd",x"48"),
   944 => (x"c2",x"c1",x"87",x"c9"),
   945 => (x"49",x"70",x"87",x"fe"),
   946 => (x"ff",x"87",x"c8",x"4a"),
   947 => (x"ff",x"c3",x"48",x"d4"),
   948 => (x"72",x"4a",x"68",x"78"),
   949 => (x"1e",x"4f",x"26",x"48"),
   950 => (x"bf",x"c0",x"df",x"c3"),
   951 => (x"05",x"a8",x"dd",x"48"),
   952 => (x"c2",x"c1",x"87",x"c6"),
   953 => (x"87",x"d9",x"87",x"ca"),
   954 => (x"c3",x"48",x"d4",x"ff"),
   955 => (x"d0",x"ff",x"78",x"ff"),
   956 => (x"78",x"e1",x"c8",x"48"),
   957 => (x"d4",x"48",x"d4",x"ff"),
   958 => (x"ff",x"de",x"c3",x"78"),
   959 => (x"bf",x"d4",x"ff",x"48"),
   960 => (x"1e",x"4f",x"26",x"50"),
   961 => (x"c0",x"48",x"d0",x"ff"),
   962 => (x"4f",x"26",x"78",x"e0"),
   963 => (x"87",x"e7",x"fe",x"1e"),
   964 => (x"02",x"99",x"49",x"70"),
   965 => (x"fb",x"c0",x"87",x"c6"),
   966 => (x"87",x"f1",x"05",x"a9"),
   967 => (x"4f",x"26",x"48",x"71"),
   968 => (x"5c",x"5b",x"5e",x"0e"),
   969 => (x"c0",x"4b",x"71",x"0e"),
   970 => (x"87",x"cb",x"fe",x"4c"),
   971 => (x"02",x"99",x"49",x"70"),
   972 => (x"c0",x"87",x"f9",x"c0"),
   973 => (x"c0",x"02",x"a9",x"ec"),
   974 => (x"fb",x"c0",x"87",x"f2"),
   975 => (x"eb",x"c0",x"02",x"a9"),
   976 => (x"b7",x"66",x"cc",x"87"),
   977 => (x"87",x"c7",x"03",x"ac"),
   978 => (x"c2",x"02",x"66",x"d0"),
   979 => (x"71",x"53",x"71",x"87"),
   980 => (x"87",x"c2",x"02",x"99"),
   981 => (x"de",x"fd",x"84",x"c1"),
   982 => (x"99",x"49",x"70",x"87"),
   983 => (x"c0",x"87",x"cd",x"02"),
   984 => (x"c7",x"02",x"a9",x"ec"),
   985 => (x"a9",x"fb",x"c0",x"87"),
   986 => (x"87",x"d5",x"ff",x"05"),
   987 => (x"c3",x"02",x"66",x"d0"),
   988 => (x"7b",x"97",x"c0",x"87"),
   989 => (x"05",x"a9",x"ec",x"c0"),
   990 => (x"4a",x"74",x"87",x"c4"),
   991 => (x"4a",x"74",x"87",x"c5"),
   992 => (x"72",x"8a",x"0a",x"c0"),
   993 => (x"26",x"87",x"c2",x"48"),
   994 => (x"26",x"4c",x"26",x"4d"),
   995 => (x"1e",x"4f",x"26",x"4b"),
   996 => (x"70",x"87",x"e4",x"fc"),
   997 => (x"b7",x"f0",x"c0",x"49"),
   998 => (x"87",x"ca",x"04",x"a9"),
   999 => (x"a9",x"b7",x"f9",x"c0"),
  1000 => (x"c0",x"87",x"c3",x"01"),
  1001 => (x"c1",x"c1",x"89",x"f0"),
  1002 => (x"ca",x"04",x"a9",x"b7"),
  1003 => (x"b7",x"da",x"c1",x"87"),
  1004 => (x"87",x"c3",x"01",x"a9"),
  1005 => (x"71",x"89",x"f7",x"c0"),
  1006 => (x"0e",x"4f",x"26",x"48"),
  1007 => (x"0e",x"5c",x"5b",x"5e"),
  1008 => (x"d4",x"ff",x"4a",x"71"),
  1009 => (x"c0",x"49",x"72",x"4c"),
  1010 => (x"4b",x"70",x"87",x"ea"),
  1011 => (x"87",x"c2",x"02",x"9b"),
  1012 => (x"d0",x"ff",x"8b",x"c1"),
  1013 => (x"78",x"c5",x"c8",x"48"),
  1014 => (x"73",x"7c",x"d5",x"c1"),
  1015 => (x"c1",x"31",x"c6",x"49"),
  1016 => (x"bf",x"97",x"e1",x"ec"),
  1017 => (x"b0",x"71",x"48",x"4a"),
  1018 => (x"d0",x"ff",x"7c",x"70"),
  1019 => (x"73",x"78",x"c4",x"48"),
  1020 => (x"87",x"d5",x"fe",x"48"),
  1021 => (x"5c",x"5b",x"5e",x"0e"),
  1022 => (x"86",x"f4",x"0e",x"5d"),
  1023 => (x"a6",x"c4",x"4c",x"71"),
  1024 => (x"c8",x"78",x"c0",x"48"),
  1025 => (x"97",x"6e",x"7e",x"a4"),
  1026 => (x"c1",x"c1",x"49",x"bf"),
  1027 => (x"87",x"dd",x"05",x"a9"),
  1028 => (x"97",x"49",x"a4",x"c9"),
  1029 => (x"d2",x"c1",x"49",x"69"),
  1030 => (x"87",x"d1",x"05",x"a9"),
  1031 => (x"97",x"49",x"a4",x"ca"),
  1032 => (x"c3",x"c1",x"49",x"69"),
  1033 => (x"87",x"c5",x"05",x"a9"),
  1034 => (x"e1",x"c2",x"48",x"df"),
  1035 => (x"87",x"e7",x"fa",x"87"),
  1036 => (x"c3",x"c1",x"4b",x"c0"),
  1037 => (x"49",x"bf",x"97",x"d3"),
  1038 => (x"cf",x"04",x"a9",x"c0"),
  1039 => (x"87",x"cc",x"fb",x"87"),
  1040 => (x"c3",x"c1",x"83",x"c1"),
  1041 => (x"49",x"bf",x"97",x"d3"),
  1042 => (x"87",x"f1",x"06",x"ab"),
  1043 => (x"97",x"d3",x"c3",x"c1"),
  1044 => (x"87",x"cf",x"02",x"bf"),
  1045 => (x"70",x"87",x"e0",x"f9"),
  1046 => (x"c6",x"02",x"99",x"49"),
  1047 => (x"a9",x"ec",x"c0",x"87"),
  1048 => (x"c0",x"87",x"f1",x"05"),
  1049 => (x"87",x"cf",x"f9",x"4b"),
  1050 => (x"ca",x"f9",x"4d",x"70"),
  1051 => (x"58",x"a6",x"cc",x"87"),
  1052 => (x"70",x"87",x"c4",x"f9"),
  1053 => (x"6e",x"83",x"c1",x"4a"),
  1054 => (x"ad",x"49",x"bf",x"97"),
  1055 => (x"c0",x"87",x"c7",x"02"),
  1056 => (x"c0",x"05",x"ad",x"ff"),
  1057 => (x"a4",x"c9",x"87",x"ea"),
  1058 => (x"49",x"69",x"97",x"49"),
  1059 => (x"02",x"a9",x"66",x"c8"),
  1060 => (x"c0",x"48",x"87",x"c7"),
  1061 => (x"d7",x"05",x"a8",x"ff"),
  1062 => (x"49",x"a4",x"ca",x"87"),
  1063 => (x"aa",x"49",x"69",x"97"),
  1064 => (x"c0",x"87",x"c6",x"02"),
  1065 => (x"c7",x"05",x"aa",x"ff"),
  1066 => (x"48",x"a6",x"c4",x"87"),
  1067 => (x"87",x"d3",x"78",x"c1"),
  1068 => (x"02",x"ad",x"ec",x"c0"),
  1069 => (x"fb",x"c0",x"87",x"c6"),
  1070 => (x"87",x"c7",x"05",x"ad"),
  1071 => (x"a6",x"c4",x"4b",x"c0"),
  1072 => (x"c4",x"78",x"c1",x"48"),
  1073 => (x"dc",x"fe",x"02",x"66"),
  1074 => (x"87",x"f7",x"f8",x"87"),
  1075 => (x"8e",x"f4",x"48",x"73"),
  1076 => (x"00",x"87",x"f4",x"fa"),
  1077 => (x"5c",x"5b",x"5e",x"0e"),
  1078 => (x"71",x"1e",x"0e",x"5d"),
  1079 => (x"4b",x"d4",x"ff",x"4d"),
  1080 => (x"df",x"c3",x"1e",x"75"),
  1081 => (x"df",x"ff",x"49",x"c4"),
  1082 => (x"86",x"c4",x"87",x"f7"),
  1083 => (x"c4",x"02",x"98",x"70"),
  1084 => (x"df",x"c3",x"87",x"cb"),
  1085 => (x"75",x"4c",x"bf",x"cc"),
  1086 => (x"87",x"ff",x"fa",x"49"),
  1087 => (x"c0",x"05",x"a8",x"de"),
  1088 => (x"49",x"75",x"87",x"eb"),
  1089 => (x"87",x"da",x"f7",x"c0"),
  1090 => (x"db",x"02",x"98",x"70"),
  1091 => (x"e8",x"e3",x"c3",x"87"),
  1092 => (x"e1",x"c0",x"1e",x"bf"),
  1093 => (x"e9",x"f4",x"c0",x"49"),
  1094 => (x"c1",x"86",x"c4",x"87"),
  1095 => (x"c0",x"48",x"e1",x"ec"),
  1096 => (x"f4",x"e3",x"c3",x"50"),
  1097 => (x"87",x"ec",x"fe",x"49"),
  1098 => (x"d2",x"c3",x"48",x"c1"),
  1099 => (x"48",x"d0",x"ff",x"87"),
  1100 => (x"c1",x"78",x"c5",x"c8"),
  1101 => (x"4a",x"c0",x"7b",x"d6"),
  1102 => (x"11",x"49",x"a2",x"75"),
  1103 => (x"cb",x"82",x"c1",x"7b"),
  1104 => (x"f3",x"04",x"aa",x"b7"),
  1105 => (x"c3",x"4a",x"cc",x"87"),
  1106 => (x"82",x"c1",x"7b",x"ff"),
  1107 => (x"aa",x"b7",x"e0",x"c0"),
  1108 => (x"ff",x"87",x"f4",x"04"),
  1109 => (x"78",x"c4",x"48",x"d0"),
  1110 => (x"c8",x"7b",x"ff",x"c3"),
  1111 => (x"d3",x"c1",x"78",x"c5"),
  1112 => (x"c4",x"7b",x"c1",x"7b"),
  1113 => (x"02",x"9c",x"74",x"78"),
  1114 => (x"c3",x"87",x"c0",x"c2"),
  1115 => (x"c8",x"7e",x"ce",x"d2"),
  1116 => (x"c0",x"8c",x"4d",x"c0"),
  1117 => (x"c6",x"03",x"ac",x"b7"),
  1118 => (x"a4",x"c0",x"c8",x"87"),
  1119 => (x"c8",x"4c",x"c0",x"4d"),
  1120 => (x"dc",x"05",x"ad",x"c0"),
  1121 => (x"ff",x"de",x"c3",x"87"),
  1122 => (x"d0",x"49",x"bf",x"97"),
  1123 => (x"87",x"d1",x"02",x"99"),
  1124 => (x"df",x"c3",x"1e",x"c0"),
  1125 => (x"dd",x"e0",x"49",x"c4"),
  1126 => (x"70",x"86",x"c4",x"87"),
  1127 => (x"ee",x"c0",x"4a",x"49"),
  1128 => (x"ce",x"d2",x"c3",x"87"),
  1129 => (x"c4",x"df",x"c3",x"1e"),
  1130 => (x"87",x"ca",x"e0",x"49"),
  1131 => (x"49",x"70",x"86",x"c4"),
  1132 => (x"48",x"d0",x"ff",x"4a"),
  1133 => (x"c1",x"78",x"c5",x"c8"),
  1134 => (x"97",x"6e",x"7b",x"d4"),
  1135 => (x"48",x"6e",x"7b",x"bf"),
  1136 => (x"7e",x"70",x"80",x"c1"),
  1137 => (x"ff",x"05",x"8d",x"c1"),
  1138 => (x"d0",x"ff",x"87",x"f0"),
  1139 => (x"72",x"78",x"c4",x"48"),
  1140 => (x"87",x"c5",x"05",x"9a"),
  1141 => (x"e6",x"c0",x"48",x"c0"),
  1142 => (x"c3",x"1e",x"c1",x"87"),
  1143 => (x"ff",x"49",x"c4",x"df"),
  1144 => (x"c4",x"87",x"f9",x"dd"),
  1145 => (x"05",x"9c",x"74",x"86"),
  1146 => (x"ff",x"87",x"c0",x"fe"),
  1147 => (x"c5",x"c8",x"48",x"d0"),
  1148 => (x"7b",x"d3",x"c1",x"78"),
  1149 => (x"78",x"c4",x"7b",x"c0"),
  1150 => (x"c2",x"c0",x"48",x"c1"),
  1151 => (x"26",x"48",x"c0",x"87"),
  1152 => (x"4c",x"26",x"4d",x"26"),
  1153 => (x"4f",x"26",x"4b",x"26"),
  1154 => (x"5c",x"5b",x"5e",x"0e"),
  1155 => (x"71",x"1e",x"0e",x"5d"),
  1156 => (x"4d",x"4c",x"c0",x"4b"),
  1157 => (x"e8",x"c0",x"04",x"ab"),
  1158 => (x"f4",x"ff",x"c0",x"87"),
  1159 => (x"02",x"9d",x"75",x"1e"),
  1160 => (x"4a",x"c0",x"87",x"c4"),
  1161 => (x"4a",x"c1",x"87",x"c2"),
  1162 => (x"d0",x"ea",x"49",x"72"),
  1163 => (x"70",x"86",x"c4",x"87"),
  1164 => (x"6e",x"84",x"c1",x"7e"),
  1165 => (x"73",x"87",x"c2",x"05"),
  1166 => (x"73",x"85",x"c1",x"4c"),
  1167 => (x"d8",x"ff",x"06",x"ac"),
  1168 => (x"26",x"48",x"6e",x"87"),
  1169 => (x"0e",x"87",x"f9",x"fe"),
  1170 => (x"0e",x"5c",x"5b",x"5e"),
  1171 => (x"66",x"cc",x"4b",x"71"),
  1172 => (x"4c",x"87",x"d8",x"02"),
  1173 => (x"02",x"8c",x"f0",x"c0"),
  1174 => (x"4a",x"74",x"87",x"d8"),
  1175 => (x"d1",x"02",x"8a",x"c1"),
  1176 => (x"cd",x"02",x"8a",x"87"),
  1177 => (x"c9",x"02",x"8a",x"87"),
  1178 => (x"73",x"87",x"d1",x"87"),
  1179 => (x"87",x"e4",x"f9",x"49"),
  1180 => (x"1e",x"74",x"87",x"ca"),
  1181 => (x"ff",x"c1",x"49",x"73"),
  1182 => (x"86",x"c4",x"87",x"e9"),
  1183 => (x"0e",x"87",x"c3",x"fe"),
  1184 => (x"5d",x"5c",x"5b",x"5e"),
  1185 => (x"4c",x"71",x"1e",x"0e"),
  1186 => (x"c3",x"91",x"de",x"49"),
  1187 => (x"71",x"4d",x"ec",x"df"),
  1188 => (x"02",x"6d",x"97",x"85"),
  1189 => (x"c3",x"87",x"dc",x"c1"),
  1190 => (x"4a",x"bf",x"d8",x"df"),
  1191 => (x"49",x"72",x"82",x"74"),
  1192 => (x"70",x"87",x"e5",x"fd"),
  1193 => (x"c0",x"02",x"6e",x"7e"),
  1194 => (x"df",x"c3",x"87",x"f2"),
  1195 => (x"4a",x"6e",x"4b",x"e0"),
  1196 => (x"f7",x"fe",x"49",x"cb"),
  1197 => (x"4b",x"74",x"87",x"f2"),
  1198 => (x"ec",x"c1",x"93",x"cb"),
  1199 => (x"83",x"c4",x"83",x"f1"),
  1200 => (x"7b",x"f7",x"cb",x"c1"),
  1201 => (x"cc",x"c1",x"49",x"74"),
  1202 => (x"7b",x"75",x"87",x"c5"),
  1203 => (x"97",x"e2",x"ec",x"c1"),
  1204 => (x"c3",x"1e",x"49",x"bf"),
  1205 => (x"fd",x"49",x"e0",x"df"),
  1206 => (x"86",x"c4",x"87",x"ed"),
  1207 => (x"cb",x"c1",x"49",x"74"),
  1208 => (x"49",x"c0",x"87",x"ed"),
  1209 => (x"87",x"cc",x"cd",x"c1"),
  1210 => (x"48",x"c0",x"df",x"c3"),
  1211 => (x"49",x"c1",x"78",x"c0"),
  1212 => (x"26",x"87",x"cf",x"dd"),
  1213 => (x"4c",x"87",x"c9",x"fc"),
  1214 => (x"69",x"64",x"61",x"6f"),
  1215 => (x"2e",x"2e",x"67",x"6e"),
  1216 => (x"5e",x"0e",x"00",x"2e"),
  1217 => (x"71",x"0e",x"5c",x"5b"),
  1218 => (x"df",x"c3",x"4a",x"4b"),
  1219 => (x"72",x"82",x"bf",x"d8"),
  1220 => (x"87",x"f4",x"fb",x"49"),
  1221 => (x"02",x"9c",x"4c",x"70"),
  1222 => (x"e5",x"49",x"87",x"c4"),
  1223 => (x"df",x"c3",x"87",x"e7"),
  1224 => (x"78",x"c0",x"48",x"d8"),
  1225 => (x"d9",x"dc",x"49",x"c1"),
  1226 => (x"87",x"d6",x"fb",x"87"),
  1227 => (x"5c",x"5b",x"5e",x"0e"),
  1228 => (x"86",x"f4",x"0e",x"5d"),
  1229 => (x"4d",x"ce",x"d2",x"c3"),
  1230 => (x"a6",x"c4",x"4c",x"c0"),
  1231 => (x"c3",x"78",x"c0",x"48"),
  1232 => (x"49",x"bf",x"d8",x"df"),
  1233 => (x"c1",x"06",x"a9",x"c0"),
  1234 => (x"d2",x"c3",x"87",x"c1"),
  1235 => (x"02",x"98",x"48",x"ce"),
  1236 => (x"c0",x"87",x"f8",x"c0"),
  1237 => (x"c8",x"1e",x"f4",x"ff"),
  1238 => (x"87",x"c7",x"02",x"66"),
  1239 => (x"c0",x"48",x"a6",x"c4"),
  1240 => (x"c4",x"87",x"c5",x"78"),
  1241 => (x"78",x"c1",x"48",x"a6"),
  1242 => (x"e5",x"49",x"66",x"c4"),
  1243 => (x"86",x"c4",x"87",x"cf"),
  1244 => (x"84",x"c1",x"4d",x"70"),
  1245 => (x"c1",x"48",x"66",x"c4"),
  1246 => (x"58",x"a6",x"c8",x"80"),
  1247 => (x"bf",x"d8",x"df",x"c3"),
  1248 => (x"c6",x"03",x"ac",x"49"),
  1249 => (x"05",x"9d",x"75",x"87"),
  1250 => (x"c0",x"87",x"c8",x"ff"),
  1251 => (x"02",x"9d",x"75",x"4c"),
  1252 => (x"c0",x"87",x"e0",x"c3"),
  1253 => (x"c8",x"1e",x"f4",x"ff"),
  1254 => (x"87",x"c7",x"02",x"66"),
  1255 => (x"c0",x"48",x"a6",x"cc"),
  1256 => (x"cc",x"87",x"c5",x"78"),
  1257 => (x"78",x"c1",x"48",x"a6"),
  1258 => (x"e4",x"49",x"66",x"cc"),
  1259 => (x"86",x"c4",x"87",x"cf"),
  1260 => (x"02",x"6e",x"7e",x"70"),
  1261 => (x"6e",x"87",x"e9",x"c2"),
  1262 => (x"97",x"81",x"cb",x"49"),
  1263 => (x"99",x"d0",x"49",x"69"),
  1264 => (x"87",x"d6",x"c1",x"02"),
  1265 => (x"4a",x"c2",x"cc",x"c1"),
  1266 => (x"91",x"cb",x"49",x"74"),
  1267 => (x"81",x"f1",x"ec",x"c1"),
  1268 => (x"81",x"c8",x"79",x"72"),
  1269 => (x"74",x"51",x"ff",x"c3"),
  1270 => (x"c3",x"91",x"de",x"49"),
  1271 => (x"71",x"4d",x"ec",x"df"),
  1272 => (x"97",x"c1",x"c2",x"85"),
  1273 => (x"49",x"a5",x"c1",x"7d"),
  1274 => (x"c3",x"51",x"e0",x"c0"),
  1275 => (x"bf",x"97",x"de",x"da"),
  1276 => (x"c1",x"87",x"d2",x"02"),
  1277 => (x"4b",x"a5",x"c2",x"84"),
  1278 => (x"4a",x"de",x"da",x"c3"),
  1279 => (x"f2",x"fe",x"49",x"db"),
  1280 => (x"db",x"c1",x"87",x"e6"),
  1281 => (x"49",x"a5",x"cd",x"87"),
  1282 => (x"84",x"c1",x"51",x"c0"),
  1283 => (x"6e",x"4b",x"a5",x"c2"),
  1284 => (x"fe",x"49",x"cb",x"4a"),
  1285 => (x"c1",x"87",x"d1",x"f2"),
  1286 => (x"c9",x"c1",x"87",x"c6"),
  1287 => (x"49",x"74",x"4a",x"ff"),
  1288 => (x"ec",x"c1",x"91",x"cb"),
  1289 => (x"79",x"72",x"81",x"f1"),
  1290 => (x"97",x"de",x"da",x"c3"),
  1291 => (x"87",x"d8",x"02",x"bf"),
  1292 => (x"91",x"de",x"49",x"74"),
  1293 => (x"df",x"c3",x"84",x"c1"),
  1294 => (x"83",x"71",x"4b",x"ec"),
  1295 => (x"4a",x"de",x"da",x"c3"),
  1296 => (x"f1",x"fe",x"49",x"dd"),
  1297 => (x"87",x"d8",x"87",x"e2"),
  1298 => (x"93",x"de",x"4b",x"74"),
  1299 => (x"83",x"ec",x"df",x"c3"),
  1300 => (x"c0",x"49",x"a3",x"cb"),
  1301 => (x"73",x"84",x"c1",x"51"),
  1302 => (x"49",x"cb",x"4a",x"6e"),
  1303 => (x"87",x"c8",x"f1",x"fe"),
  1304 => (x"c1",x"48",x"66",x"c4"),
  1305 => (x"58",x"a6",x"c8",x"80"),
  1306 => (x"c0",x"03",x"ac",x"c7"),
  1307 => (x"05",x"6e",x"87",x"c5"),
  1308 => (x"74",x"87",x"e0",x"fc"),
  1309 => (x"f6",x"8e",x"f4",x"48"),
  1310 => (x"73",x"1e",x"87",x"c6"),
  1311 => (x"49",x"4b",x"71",x"1e"),
  1312 => (x"ec",x"c1",x"91",x"cb"),
  1313 => (x"a1",x"c8",x"81",x"f1"),
  1314 => (x"e1",x"ec",x"c1",x"4a"),
  1315 => (x"c9",x"50",x"12",x"48"),
  1316 => (x"c3",x"c1",x"4a",x"a1"),
  1317 => (x"50",x"12",x"48",x"d3"),
  1318 => (x"ec",x"c1",x"81",x"ca"),
  1319 => (x"50",x"11",x"48",x"e2"),
  1320 => (x"97",x"e2",x"ec",x"c1"),
  1321 => (x"c0",x"1e",x"49",x"bf"),
  1322 => (x"87",x"db",x"f6",x"49"),
  1323 => (x"48",x"c0",x"df",x"c3"),
  1324 => (x"49",x"c1",x"78",x"de"),
  1325 => (x"26",x"87",x"cb",x"d6"),
  1326 => (x"1e",x"87",x"c9",x"f5"),
  1327 => (x"cb",x"49",x"4a",x"71"),
  1328 => (x"f1",x"ec",x"c1",x"91"),
  1329 => (x"11",x"81",x"c8",x"81"),
  1330 => (x"c4",x"df",x"c3",x"48"),
  1331 => (x"d8",x"df",x"c3",x"58"),
  1332 => (x"c1",x"78",x"c0",x"48"),
  1333 => (x"87",x"ea",x"d5",x"49"),
  1334 => (x"c0",x"1e",x"4f",x"26"),
  1335 => (x"d3",x"c5",x"c1",x"49"),
  1336 => (x"1e",x"4f",x"26",x"87"),
  1337 => (x"d2",x"02",x"99",x"71"),
  1338 => (x"c6",x"ee",x"c1",x"87"),
  1339 => (x"f7",x"50",x"c0",x"48"),
  1340 => (x"fb",x"d2",x"c1",x"80"),
  1341 => (x"ea",x"ec",x"c1",x"40"),
  1342 => (x"c1",x"87",x"ce",x"78"),
  1343 => (x"c1",x"48",x"c2",x"ee"),
  1344 => (x"fc",x"78",x"e3",x"ec"),
  1345 => (x"da",x"d3",x"c1",x"80"),
  1346 => (x"0e",x"4f",x"26",x"78"),
  1347 => (x"0e",x"5c",x"5b",x"5e"),
  1348 => (x"cb",x"4a",x"4c",x"71"),
  1349 => (x"f1",x"ec",x"c1",x"92"),
  1350 => (x"49",x"a2",x"c8",x"82"),
  1351 => (x"97",x"4b",x"a2",x"c9"),
  1352 => (x"97",x"1e",x"4b",x"6b"),
  1353 => (x"ca",x"1e",x"49",x"69"),
  1354 => (x"c0",x"49",x"12",x"82"),
  1355 => (x"c0",x"87",x"f3",x"e5"),
  1356 => (x"87",x"ce",x"d4",x"49"),
  1357 => (x"c2",x"c1",x"49",x"74"),
  1358 => (x"8e",x"f8",x"87",x"d5"),
  1359 => (x"1e",x"87",x"c3",x"f3"),
  1360 => (x"4b",x"71",x"1e",x"73"),
  1361 => (x"87",x"c3",x"ff",x"49"),
  1362 => (x"fe",x"fe",x"49",x"73"),
  1363 => (x"87",x"f4",x"f2",x"87"),
  1364 => (x"71",x"1e",x"73",x"1e"),
  1365 => (x"4a",x"a3",x"c6",x"4b"),
  1366 => (x"c1",x"87",x"db",x"02"),
  1367 => (x"87",x"d6",x"02",x"8a"),
  1368 => (x"da",x"c1",x"02",x"8a"),
  1369 => (x"c0",x"02",x"8a",x"87"),
  1370 => (x"02",x"8a",x"87",x"fc"),
  1371 => (x"8a",x"87",x"e1",x"c0"),
  1372 => (x"c1",x"87",x"cb",x"02"),
  1373 => (x"49",x"c7",x"87",x"db"),
  1374 => (x"c1",x"87",x"c0",x"fd"),
  1375 => (x"df",x"c3",x"87",x"de"),
  1376 => (x"c1",x"02",x"bf",x"d8"),
  1377 => (x"c1",x"48",x"87",x"cb"),
  1378 => (x"dc",x"df",x"c3",x"88"),
  1379 => (x"87",x"c1",x"c1",x"58"),
  1380 => (x"bf",x"dc",x"df",x"c3"),
  1381 => (x"87",x"f9",x"c0",x"02"),
  1382 => (x"bf",x"d8",x"df",x"c3"),
  1383 => (x"c3",x"80",x"c1",x"48"),
  1384 => (x"c0",x"58",x"dc",x"df"),
  1385 => (x"df",x"c3",x"87",x"eb"),
  1386 => (x"c6",x"49",x"bf",x"d8"),
  1387 => (x"dc",x"df",x"c3",x"89"),
  1388 => (x"a9",x"b7",x"c0",x"59"),
  1389 => (x"c3",x"87",x"da",x"03"),
  1390 => (x"c0",x"48",x"d8",x"df"),
  1391 => (x"c3",x"87",x"d2",x"78"),
  1392 => (x"02",x"bf",x"dc",x"df"),
  1393 => (x"df",x"c3",x"87",x"cb"),
  1394 => (x"c6",x"48",x"bf",x"d8"),
  1395 => (x"dc",x"df",x"c3",x"80"),
  1396 => (x"d1",x"49",x"c0",x"58"),
  1397 => (x"49",x"73",x"87",x"ec"),
  1398 => (x"87",x"f3",x"ff",x"c0"),
  1399 => (x"1e",x"87",x"e5",x"f0"),
  1400 => (x"4b",x"71",x"1e",x"73"),
  1401 => (x"48",x"c0",x"df",x"c3"),
  1402 => (x"49",x"c0",x"78",x"dd"),
  1403 => (x"73",x"87",x"d3",x"d1"),
  1404 => (x"da",x"ff",x"c0",x"49"),
  1405 => (x"87",x"cc",x"f0",x"87"),
  1406 => (x"5c",x"5b",x"5e",x"0e"),
  1407 => (x"cc",x"4c",x"71",x"0e"),
  1408 => (x"4b",x"74",x"1e",x"66"),
  1409 => (x"ec",x"c1",x"93",x"cb"),
  1410 => (x"a3",x"c4",x"83",x"f1"),
  1411 => (x"fe",x"49",x"6a",x"4a"),
  1412 => (x"c1",x"87",x"e5",x"ea"),
  1413 => (x"c8",x"7b",x"fa",x"d1"),
  1414 => (x"66",x"d4",x"49",x"a3"),
  1415 => (x"49",x"a3",x"c9",x"51"),
  1416 => (x"ca",x"51",x"66",x"d8"),
  1417 => (x"66",x"dc",x"49",x"a3"),
  1418 => (x"d5",x"ef",x"26",x"51"),
  1419 => (x"5b",x"5e",x"0e",x"87"),
  1420 => (x"ff",x"0e",x"5d",x"5c"),
  1421 => (x"a6",x"dc",x"86",x"cc"),
  1422 => (x"48",x"a6",x"c8",x"59"),
  1423 => (x"80",x"c4",x"78",x"c0"),
  1424 => (x"78",x"66",x"c8",x"c1"),
  1425 => (x"78",x"c1",x"80",x"c4"),
  1426 => (x"78",x"c1",x"80",x"c4"),
  1427 => (x"48",x"dc",x"df",x"c3"),
  1428 => (x"df",x"c3",x"78",x"c1"),
  1429 => (x"de",x"48",x"bf",x"c0"),
  1430 => (x"87",x"cb",x"05",x"a8"),
  1431 => (x"70",x"87",x"cd",x"f3"),
  1432 => (x"59",x"a6",x"cc",x"49"),
  1433 => (x"e1",x"87",x"d6",x"ce"),
  1434 => (x"df",x"e2",x"87",x"ed"),
  1435 => (x"87",x"c7",x"e1",x"87"),
  1436 => (x"fb",x"c0",x"4c",x"70"),
  1437 => (x"d8",x"c1",x"02",x"ac"),
  1438 => (x"05",x"66",x"d8",x"87"),
  1439 => (x"c0",x"87",x"ca",x"c1"),
  1440 => (x"1e",x"c1",x"1e",x"1e"),
  1441 => (x"1e",x"e4",x"ee",x"c1"),
  1442 => (x"eb",x"fd",x"49",x"c0"),
  1443 => (x"c0",x"86",x"d0",x"87"),
  1444 => (x"d9",x"02",x"ac",x"fb"),
  1445 => (x"66",x"c4",x"c1",x"87"),
  1446 => (x"6a",x"82",x"c4",x"4a"),
  1447 => (x"74",x"81",x"c7",x"49"),
  1448 => (x"d8",x"1e",x"c1",x"51"),
  1449 => (x"c8",x"49",x"6a",x"1e"),
  1450 => (x"87",x"f4",x"e1",x"81"),
  1451 => (x"c8",x"c1",x"86",x"c8"),
  1452 => (x"a8",x"c0",x"48",x"66"),
  1453 => (x"c8",x"87",x"c7",x"01"),
  1454 => (x"78",x"c1",x"48",x"a6"),
  1455 => (x"c8",x"c1",x"87",x"ce"),
  1456 => (x"88",x"c1",x"48",x"66"),
  1457 => (x"c3",x"58",x"a6",x"d0"),
  1458 => (x"87",x"c0",x"e1",x"87"),
  1459 => (x"c2",x"48",x"a6",x"d0"),
  1460 => (x"02",x"9c",x"74",x"78"),
  1461 => (x"c8",x"87",x"e2",x"cc"),
  1462 => (x"cc",x"c1",x"48",x"66"),
  1463 => (x"cc",x"03",x"a8",x"66"),
  1464 => (x"a6",x"c4",x"87",x"d7"),
  1465 => (x"d8",x"78",x"c0",x"48"),
  1466 => (x"ff",x"78",x"c0",x"80"),
  1467 => (x"70",x"87",x"c8",x"df"),
  1468 => (x"48",x"66",x"d8",x"4c"),
  1469 => (x"c6",x"05",x"a8",x"dd"),
  1470 => (x"48",x"a6",x"dc",x"87"),
  1471 => (x"c1",x"78",x"66",x"d8"),
  1472 => (x"c0",x"05",x"ac",x"d0"),
  1473 => (x"de",x"ff",x"87",x"eb"),
  1474 => (x"de",x"ff",x"87",x"ed"),
  1475 => (x"4c",x"70",x"87",x"e9"),
  1476 => (x"05",x"ac",x"ec",x"c0"),
  1477 => (x"df",x"ff",x"87",x"c6"),
  1478 => (x"4c",x"70",x"87",x"f2"),
  1479 => (x"05",x"ac",x"d0",x"c1"),
  1480 => (x"66",x"d4",x"87",x"c8"),
  1481 => (x"d8",x"80",x"c1",x"48"),
  1482 => (x"d0",x"c1",x"58",x"a6"),
  1483 => (x"d5",x"ff",x"02",x"ac"),
  1484 => (x"a6",x"e0",x"c0",x"87"),
  1485 => (x"78",x"66",x"d8",x"48"),
  1486 => (x"c0",x"48",x"66",x"dc"),
  1487 => (x"05",x"a8",x"66",x"e0"),
  1488 => (x"c0",x"87",x"c8",x"ca"),
  1489 => (x"c0",x"48",x"a6",x"e4"),
  1490 => (x"c0",x"80",x"c4",x"78"),
  1491 => (x"c0",x"4d",x"74",x"78"),
  1492 => (x"c9",x"02",x"8d",x"fb"),
  1493 => (x"8d",x"c9",x"87",x"ce"),
  1494 => (x"c2",x"87",x"db",x"02"),
  1495 => (x"f7",x"c1",x"02",x"8d"),
  1496 => (x"02",x"8d",x"c9",x"87"),
  1497 => (x"c4",x"87",x"d1",x"c4"),
  1498 => (x"c2",x"c1",x"02",x"8d"),
  1499 => (x"02",x"8d",x"c1",x"87"),
  1500 => (x"c8",x"87",x"c5",x"c4"),
  1501 => (x"66",x"c8",x"87",x"e8"),
  1502 => (x"c1",x"91",x"cb",x"49"),
  1503 => (x"c4",x"81",x"66",x"c4"),
  1504 => (x"7e",x"6a",x"4a",x"a1"),
  1505 => (x"e8",x"c1",x"1e",x"71"),
  1506 => (x"66",x"c4",x"48",x"f5"),
  1507 => (x"4a",x"a1",x"cc",x"49"),
  1508 => (x"aa",x"71",x"41",x"20"),
  1509 => (x"87",x"f8",x"ff",x"05"),
  1510 => (x"49",x"26",x"51",x"10"),
  1511 => (x"79",x"df",x"d7",x"c1"),
  1512 => (x"87",x"e8",x"dd",x"ff"),
  1513 => (x"e8",x"c0",x"4c",x"70"),
  1514 => (x"78",x"c1",x"48",x"a6"),
  1515 => (x"c4",x"87",x"f5",x"c7"),
  1516 => (x"f0",x"c0",x"48",x"a6"),
  1517 => (x"fe",x"db",x"ff",x"78"),
  1518 => (x"c0",x"4c",x"70",x"87"),
  1519 => (x"c0",x"02",x"ac",x"ec"),
  1520 => (x"a6",x"c8",x"87",x"c3"),
  1521 => (x"ac",x"ec",x"c0",x"5c"),
  1522 => (x"ff",x"87",x"cd",x"02"),
  1523 => (x"70",x"87",x"e8",x"db"),
  1524 => (x"ac",x"ec",x"c0",x"4c"),
  1525 => (x"87",x"f3",x"ff",x"05"),
  1526 => (x"02",x"ac",x"ec",x"c0"),
  1527 => (x"ff",x"87",x"c4",x"c0"),
  1528 => (x"c4",x"87",x"d4",x"db"),
  1529 => (x"66",x"d8",x"1e",x"66"),
  1530 => (x"66",x"d8",x"1e",x"49"),
  1531 => (x"ee",x"c1",x"1e",x"49"),
  1532 => (x"66",x"d8",x"1e",x"e4"),
  1533 => (x"87",x"c0",x"f8",x"49"),
  1534 => (x"1e",x"ca",x"1e",x"c0"),
  1535 => (x"49",x"66",x"e0",x"c0"),
  1536 => (x"dc",x"c1",x"91",x"cb"),
  1537 => (x"a6",x"d8",x"81",x"66"),
  1538 => (x"78",x"a1",x"c4",x"48"),
  1539 => (x"49",x"bf",x"66",x"d8"),
  1540 => (x"87",x"cc",x"dc",x"ff"),
  1541 => (x"b7",x"c0",x"86",x"d8"),
  1542 => (x"cb",x"c1",x"06",x"a8"),
  1543 => (x"de",x"1e",x"c1",x"87"),
  1544 => (x"bf",x"66",x"c8",x"1e"),
  1545 => (x"f7",x"db",x"ff",x"49"),
  1546 => (x"70",x"86",x"c8",x"87"),
  1547 => (x"08",x"c0",x"48",x"49"),
  1548 => (x"a6",x"ec",x"c0",x"88"),
  1549 => (x"a8",x"b7",x"c0",x"58"),
  1550 => (x"87",x"ec",x"c0",x"06"),
  1551 => (x"48",x"66",x"e8",x"c0"),
  1552 => (x"03",x"a8",x"b7",x"dd"),
  1553 => (x"6e",x"87",x"e1",x"c0"),
  1554 => (x"e8",x"c0",x"49",x"bf"),
  1555 => (x"e0",x"c0",x"81",x"66"),
  1556 => (x"66",x"e8",x"c0",x"51"),
  1557 => (x"6e",x"81",x"c1",x"49"),
  1558 => (x"c1",x"c2",x"81",x"bf"),
  1559 => (x"66",x"e8",x"c0",x"51"),
  1560 => (x"6e",x"81",x"c2",x"49"),
  1561 => (x"51",x"c0",x"81",x"bf"),
  1562 => (x"c1",x"48",x"66",x"d0"),
  1563 => (x"58",x"a6",x"d4",x"80"),
  1564 => (x"c1",x"80",x"d8",x"48"),
  1565 => (x"87",x"ec",x"c4",x"78"),
  1566 => (x"87",x"d3",x"dc",x"ff"),
  1567 => (x"58",x"a6",x"ec",x"c0"),
  1568 => (x"87",x"cb",x"dc",x"ff"),
  1569 => (x"58",x"a6",x"f0",x"c0"),
  1570 => (x"05",x"a8",x"ec",x"c0"),
  1571 => (x"a6",x"87",x"c9",x"c0"),
  1572 => (x"66",x"e8",x"c0",x"48"),
  1573 => (x"87",x"c4",x"c0",x"78"),
  1574 => (x"87",x"db",x"d8",x"ff"),
  1575 => (x"cb",x"49",x"66",x"c8"),
  1576 => (x"66",x"c4",x"c1",x"91"),
  1577 => (x"c8",x"80",x"71",x"48"),
  1578 => (x"66",x"c4",x"58",x"a6"),
  1579 => (x"c4",x"82",x"c8",x"4a"),
  1580 => (x"81",x"ca",x"49",x"66"),
  1581 => (x"51",x"66",x"e8",x"c0"),
  1582 => (x"49",x"66",x"ec",x"c0"),
  1583 => (x"e8",x"c0",x"81",x"c1"),
  1584 => (x"48",x"c1",x"89",x"66"),
  1585 => (x"49",x"70",x"30",x"71"),
  1586 => (x"97",x"71",x"89",x"c1"),
  1587 => (x"c8",x"e3",x"c3",x"7a"),
  1588 => (x"e8",x"c0",x"49",x"bf"),
  1589 => (x"6a",x"97",x"29",x"66"),
  1590 => (x"98",x"71",x"48",x"4a"),
  1591 => (x"58",x"a6",x"f4",x"c0"),
  1592 => (x"c4",x"49",x"66",x"c4"),
  1593 => (x"c0",x"7e",x"69",x"81"),
  1594 => (x"dc",x"48",x"66",x"e0"),
  1595 => (x"c0",x"02",x"a8",x"66"),
  1596 => (x"a6",x"dc",x"87",x"c8"),
  1597 => (x"c0",x"78",x"c0",x"48"),
  1598 => (x"a6",x"dc",x"87",x"c5"),
  1599 => (x"dc",x"78",x"c1",x"48"),
  1600 => (x"e0",x"c0",x"1e",x"66"),
  1601 => (x"49",x"66",x"c8",x"1e"),
  1602 => (x"87",x"d4",x"d8",x"ff"),
  1603 => (x"4c",x"70",x"86",x"c8"),
  1604 => (x"06",x"ac",x"b7",x"c0"),
  1605 => (x"6e",x"87",x"d6",x"c1"),
  1606 => (x"70",x"80",x"74",x"48"),
  1607 => (x"49",x"e0",x"c0",x"7e"),
  1608 => (x"4b",x"6e",x"89",x"74"),
  1609 => (x"4a",x"f2",x"e8",x"c1"),
  1610 => (x"fb",x"dd",x"fe",x"71"),
  1611 => (x"c2",x"48",x"6e",x"87"),
  1612 => (x"c0",x"7e",x"70",x"80"),
  1613 => (x"c1",x"48",x"66",x"e4"),
  1614 => (x"a6",x"e8",x"c0",x"80"),
  1615 => (x"66",x"f0",x"c0",x"58"),
  1616 => (x"70",x"81",x"c1",x"49"),
  1617 => (x"c5",x"c0",x"02",x"a9"),
  1618 => (x"c0",x"4d",x"c0",x"87"),
  1619 => (x"4d",x"c1",x"87",x"c2"),
  1620 => (x"a4",x"c2",x"1e",x"75"),
  1621 => (x"48",x"e0",x"c0",x"49"),
  1622 => (x"49",x"70",x"88",x"71"),
  1623 => (x"49",x"66",x"c8",x"1e"),
  1624 => (x"87",x"fc",x"d6",x"ff"),
  1625 => (x"b7",x"c0",x"86",x"c8"),
  1626 => (x"c6",x"ff",x"01",x"a8"),
  1627 => (x"66",x"e4",x"c0",x"87"),
  1628 => (x"87",x"d3",x"c0",x"02"),
  1629 => (x"c9",x"49",x"66",x"c4"),
  1630 => (x"66",x"e4",x"c0",x"81"),
  1631 => (x"48",x"66",x"c4",x"51"),
  1632 => (x"78",x"cb",x"d4",x"c1"),
  1633 => (x"c4",x"87",x"ce",x"c0"),
  1634 => (x"81",x"c9",x"49",x"66"),
  1635 => (x"66",x"c4",x"51",x"c2"),
  1636 => (x"ff",x"d4",x"c1",x"48"),
  1637 => (x"a6",x"e8",x"c0",x"78"),
  1638 => (x"c0",x"78",x"c1",x"48"),
  1639 => (x"d5",x"ff",x"87",x"c6"),
  1640 => (x"4c",x"70",x"87",x"ea"),
  1641 => (x"02",x"66",x"e8",x"c0"),
  1642 => (x"c8",x"87",x"f5",x"c0"),
  1643 => (x"66",x"cc",x"48",x"66"),
  1644 => (x"cb",x"c0",x"04",x"a8"),
  1645 => (x"48",x"66",x"c8",x"87"),
  1646 => (x"a6",x"cc",x"80",x"c1"),
  1647 => (x"87",x"e0",x"c0",x"58"),
  1648 => (x"c1",x"48",x"66",x"cc"),
  1649 => (x"58",x"a6",x"d0",x"88"),
  1650 => (x"c1",x"87",x"d5",x"c0"),
  1651 => (x"c0",x"05",x"ac",x"c6"),
  1652 => (x"66",x"d0",x"87",x"c8"),
  1653 => (x"d4",x"80",x"c1",x"48"),
  1654 => (x"d4",x"ff",x"58",x"a6"),
  1655 => (x"4c",x"70",x"87",x"ee"),
  1656 => (x"c1",x"48",x"66",x"d4"),
  1657 => (x"58",x"a6",x"d8",x"80"),
  1658 => (x"c0",x"02",x"9c",x"74"),
  1659 => (x"66",x"c8",x"87",x"cb"),
  1660 => (x"66",x"cc",x"c1",x"48"),
  1661 => (x"e9",x"f3",x"04",x"a8"),
  1662 => (x"c6",x"d4",x"ff",x"87"),
  1663 => (x"48",x"66",x"c8",x"87"),
  1664 => (x"c0",x"03",x"a8",x"c7"),
  1665 => (x"df",x"c3",x"87",x"e5"),
  1666 => (x"78",x"c0",x"48",x"dc"),
  1667 => (x"cb",x"49",x"66",x"c8"),
  1668 => (x"66",x"c4",x"c1",x"91"),
  1669 => (x"4a",x"a1",x"c4",x"81"),
  1670 => (x"52",x"c0",x"4a",x"6a"),
  1671 => (x"48",x"66",x"c8",x"79"),
  1672 => (x"a6",x"cc",x"80",x"c1"),
  1673 => (x"04",x"a8",x"c7",x"58"),
  1674 => (x"ff",x"87",x"db",x"ff"),
  1675 => (x"df",x"ff",x"8e",x"cc"),
  1676 => (x"20",x"3a",x"87",x"ce"),
  1677 => (x"50",x"49",x"44",x"00"),
  1678 => (x"69",x"77",x"53",x"20"),
  1679 => (x"65",x"68",x"63",x"74"),
  1680 => (x"73",x"1e",x"00",x"73"),
  1681 => (x"9b",x"4b",x"71",x"1e"),
  1682 => (x"c3",x"87",x"c6",x"02"),
  1683 => (x"c0",x"48",x"d8",x"df"),
  1684 => (x"c3",x"1e",x"c7",x"78"),
  1685 => (x"49",x"bf",x"d8",x"df"),
  1686 => (x"f1",x"ec",x"c1",x"1e"),
  1687 => (x"c0",x"df",x"c3",x"1e"),
  1688 => (x"c8",x"ef",x"49",x"bf"),
  1689 => (x"c3",x"86",x"cc",x"87"),
  1690 => (x"49",x"bf",x"c0",x"df"),
  1691 => (x"73",x"87",x"f4",x"e9"),
  1692 => (x"87",x"c8",x"02",x"9b"),
  1693 => (x"49",x"f1",x"ec",x"c1"),
  1694 => (x"87",x"e5",x"ee",x"c0"),
  1695 => (x"87",x"c4",x"de",x"ff"),
  1696 => (x"e1",x"ec",x"c1",x"1e"),
  1697 => (x"c1",x"50",x"c0",x"48"),
  1698 => (x"49",x"bf",x"d4",x"ee"),
  1699 => (x"87",x"c4",x"d9",x"ff"),
  1700 => (x"4f",x"26",x"48",x"c0"),
  1701 => (x"87",x"eb",x"c7",x"1e"),
  1702 => (x"e5",x"fe",x"49",x"c1"),
  1703 => (x"ee",x"e2",x"fe",x"87"),
  1704 => (x"02",x"98",x"70",x"87"),
  1705 => (x"eb",x"fe",x"87",x"cd"),
  1706 => (x"98",x"70",x"87",x"e9"),
  1707 => (x"c1",x"87",x"c4",x"02"),
  1708 => (x"c0",x"87",x"c2",x"4a"),
  1709 => (x"05",x"9a",x"72",x"4a"),
  1710 => (x"1e",x"c0",x"87",x"ce"),
  1711 => (x"49",x"e8",x"eb",x"c1"),
  1712 => (x"87",x"fe",x"f9",x"c0"),
  1713 => (x"87",x"fe",x"86",x"c4"),
  1714 => (x"87",x"f0",x"e5",x"c1"),
  1715 => (x"eb",x"c1",x"1e",x"c0"),
  1716 => (x"f9",x"c0",x"49",x"f3"),
  1717 => (x"1e",x"c0",x"87",x"ec"),
  1718 => (x"70",x"87",x"e5",x"fe"),
  1719 => (x"e1",x"f9",x"c0",x"49"),
  1720 => (x"87",x"de",x"c3",x"87"),
  1721 => (x"4f",x"26",x"8e",x"f8"),
  1722 => (x"66",x"20",x"44",x"53"),
  1723 => (x"65",x"6c",x"69",x"61"),
  1724 => (x"42",x"00",x"2e",x"64"),
  1725 => (x"69",x"74",x"6f",x"6f"),
  1726 => (x"2e",x"2e",x"67",x"6e"),
  1727 => (x"c0",x"1e",x"00",x"2e"),
  1728 => (x"c1",x"87",x"ff",x"f0"),
  1729 => (x"f6",x"87",x"c6",x"de"),
  1730 => (x"1e",x"4f",x"26",x"87"),
  1731 => (x"48",x"d8",x"df",x"c3"),
  1732 => (x"df",x"c3",x"78",x"c0"),
  1733 => (x"78",x"c0",x"48",x"c0"),
  1734 => (x"e1",x"87",x"f9",x"fd"),
  1735 => (x"26",x"48",x"c0",x"87"),
  1736 => (x"80",x"00",x"00",x"4f"),
  1737 => (x"69",x"78",x"45",x"20"),
  1738 => (x"20",x"80",x"00",x"74"),
  1739 => (x"6b",x"63",x"61",x"42"),
  1740 => (x"00",x"14",x"bb",x"00"),
  1741 => (x"00",x"37",x"ec",x"00"),
  1742 => (x"00",x"00",x"00",x"00"),
  1743 => (x"00",x"00",x"14",x"bb"),
  1744 => (x"00",x"00",x"38",x"0a"),
  1745 => (x"bb",x"00",x"00",x"00"),
  1746 => (x"28",x"00",x"00",x"14"),
  1747 => (x"00",x"00",x"00",x"38"),
  1748 => (x"14",x"bb",x"00",x"00"),
  1749 => (x"38",x"46",x"00",x"00"),
  1750 => (x"00",x"00",x"00",x"00"),
  1751 => (x"00",x"14",x"bb",x"00"),
  1752 => (x"00",x"38",x"64",x"00"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"00",x"00",x"14",x"bb"),
  1755 => (x"00",x"00",x"38",x"82"),
  1756 => (x"bb",x"00",x"00",x"00"),
  1757 => (x"a0",x"00",x"00",x"14"),
  1758 => (x"00",x"00",x"00",x"38"),
  1759 => (x"14",x"bb",x"00",x"00"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"15",x"50",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"1b",x"98"),
  1766 => (x"54",x"4f",x"4f",x"42"),
  1767 => (x"20",x"20",x"20",x"20"),
  1768 => (x"00",x"4d",x"4f",x"52"),
  1769 => (x"64",x"61",x"6f",x"4c"),
  1770 => (x"00",x"2e",x"2a",x"20"),
  1771 => (x"48",x"f0",x"fe",x"1e"),
  1772 => (x"09",x"cd",x"78",x"c0"),
  1773 => (x"4f",x"26",x"09",x"79"),
  1774 => (x"f0",x"fe",x"1e",x"1e"),
  1775 => (x"26",x"48",x"7e",x"bf"),
  1776 => (x"fe",x"1e",x"4f",x"26"),
  1777 => (x"78",x"c1",x"48",x"f0"),
  1778 => (x"fe",x"1e",x"4f",x"26"),
  1779 => (x"78",x"c0",x"48",x"f0"),
  1780 => (x"71",x"1e",x"4f",x"26"),
  1781 => (x"52",x"52",x"c0",x"4a"),
  1782 => (x"5e",x"0e",x"4f",x"26"),
  1783 => (x"0e",x"5d",x"5c",x"5b"),
  1784 => (x"4d",x"71",x"86",x"f4"),
  1785 => (x"c1",x"7e",x"6d",x"97"),
  1786 => (x"6c",x"97",x"4c",x"a5"),
  1787 => (x"58",x"a6",x"c8",x"48"),
  1788 => (x"66",x"c4",x"48",x"6e"),
  1789 => (x"87",x"c5",x"05",x"a8"),
  1790 => (x"e6",x"c0",x"48",x"ff"),
  1791 => (x"87",x"ca",x"ff",x"87"),
  1792 => (x"97",x"49",x"a5",x"c2"),
  1793 => (x"a3",x"71",x"4b",x"6c"),
  1794 => (x"4b",x"6b",x"97",x"4b"),
  1795 => (x"6e",x"7e",x"6c",x"97"),
  1796 => (x"c8",x"80",x"c1",x"48"),
  1797 => (x"98",x"c7",x"58",x"a6"),
  1798 => (x"70",x"58",x"a6",x"cc"),
  1799 => (x"e1",x"fe",x"7c",x"97"),
  1800 => (x"f4",x"48",x"73",x"87"),
  1801 => (x"26",x"4d",x"26",x"8e"),
  1802 => (x"26",x"4b",x"26",x"4c"),
  1803 => (x"5b",x"5e",x"0e",x"4f"),
  1804 => (x"86",x"f4",x"0e",x"5c"),
  1805 => (x"66",x"d8",x"4c",x"71"),
  1806 => (x"9a",x"ff",x"c3",x"4a"),
  1807 => (x"97",x"4b",x"a4",x"c2"),
  1808 => (x"a1",x"73",x"49",x"6c"),
  1809 => (x"97",x"51",x"72",x"49"),
  1810 => (x"48",x"6e",x"7e",x"6c"),
  1811 => (x"a6",x"c8",x"80",x"c1"),
  1812 => (x"cc",x"98",x"c7",x"58"),
  1813 => (x"54",x"70",x"58",x"a6"),
  1814 => (x"ca",x"ff",x"8e",x"f4"),
  1815 => (x"fd",x"1e",x"1e",x"87"),
  1816 => (x"bf",x"e0",x"87",x"e8"),
  1817 => (x"e0",x"c0",x"49",x"4a"),
  1818 => (x"cb",x"02",x"99",x"c0"),
  1819 => (x"c3",x"1e",x"72",x"87"),
  1820 => (x"fe",x"49",x"fe",x"e2"),
  1821 => (x"86",x"c4",x"87",x"f7"),
  1822 => (x"70",x"87",x"fd",x"fc"),
  1823 => (x"87",x"c2",x"fd",x"7e"),
  1824 => (x"1e",x"4f",x"26",x"26"),
  1825 => (x"49",x"fe",x"e2",x"c3"),
  1826 => (x"c1",x"87",x"c7",x"fd"),
  1827 => (x"fc",x"49",x"dd",x"f1"),
  1828 => (x"c8",x"c4",x"87",x"da"),
  1829 => (x"1e",x"4f",x"26",x"87"),
  1830 => (x"c8",x"48",x"d0",x"ff"),
  1831 => (x"d4",x"ff",x"78",x"e1"),
  1832 => (x"c4",x"78",x"c5",x"48"),
  1833 => (x"87",x"c3",x"02",x"66"),
  1834 => (x"c8",x"78",x"e0",x"c3"),
  1835 => (x"87",x"c6",x"02",x"66"),
  1836 => (x"c3",x"48",x"d4",x"ff"),
  1837 => (x"d4",x"ff",x"78",x"f0"),
  1838 => (x"ff",x"78",x"71",x"48"),
  1839 => (x"e1",x"c8",x"48",x"d0"),
  1840 => (x"78",x"e0",x"c0",x"78"),
  1841 => (x"5e",x"0e",x"4f",x"26"),
  1842 => (x"71",x"0e",x"5c",x"5b"),
  1843 => (x"fe",x"e2",x"c3",x"4c"),
  1844 => (x"87",x"c6",x"fc",x"49"),
  1845 => (x"b7",x"c0",x"4a",x"70"),
  1846 => (x"e3",x"c2",x"04",x"aa"),
  1847 => (x"aa",x"e0",x"c3",x"87"),
  1848 => (x"c1",x"87",x"c9",x"05"),
  1849 => (x"c1",x"48",x"d0",x"f6"),
  1850 => (x"87",x"d4",x"c2",x"78"),
  1851 => (x"05",x"aa",x"f0",x"c3"),
  1852 => (x"f6",x"c1",x"87",x"c9"),
  1853 => (x"78",x"c1",x"48",x"cc"),
  1854 => (x"c1",x"87",x"f5",x"c1"),
  1855 => (x"02",x"bf",x"d0",x"f6"),
  1856 => (x"4b",x"72",x"87",x"c7"),
  1857 => (x"c2",x"b3",x"c0",x"c2"),
  1858 => (x"74",x"4b",x"72",x"87"),
  1859 => (x"87",x"d1",x"05",x"9c"),
  1860 => (x"bf",x"cc",x"f6",x"c1"),
  1861 => (x"d0",x"f6",x"c1",x"1e"),
  1862 => (x"49",x"72",x"1e",x"bf"),
  1863 => (x"c8",x"87",x"f8",x"fd"),
  1864 => (x"cc",x"f6",x"c1",x"86"),
  1865 => (x"e0",x"c0",x"02",x"bf"),
  1866 => (x"c4",x"49",x"73",x"87"),
  1867 => (x"c1",x"91",x"29",x"b7"),
  1868 => (x"73",x"81",x"ec",x"f7"),
  1869 => (x"c2",x"9a",x"cf",x"4a"),
  1870 => (x"72",x"48",x"c1",x"92"),
  1871 => (x"ff",x"4a",x"70",x"30"),
  1872 => (x"69",x"48",x"72",x"ba"),
  1873 => (x"db",x"79",x"70",x"98"),
  1874 => (x"c4",x"49",x"73",x"87"),
  1875 => (x"c1",x"91",x"29",x"b7"),
  1876 => (x"73",x"81",x"ec",x"f7"),
  1877 => (x"c2",x"9a",x"cf",x"4a"),
  1878 => (x"72",x"48",x"c3",x"92"),
  1879 => (x"48",x"4a",x"70",x"30"),
  1880 => (x"79",x"70",x"b0",x"69"),
  1881 => (x"48",x"d0",x"f6",x"c1"),
  1882 => (x"f6",x"c1",x"78",x"c0"),
  1883 => (x"78",x"c0",x"48",x"cc"),
  1884 => (x"49",x"fe",x"e2",x"c3"),
  1885 => (x"70",x"87",x"e3",x"f9"),
  1886 => (x"aa",x"b7",x"c0",x"4a"),
  1887 => (x"87",x"dd",x"fd",x"03"),
  1888 => (x"87",x"c2",x"48",x"c0"),
  1889 => (x"4c",x"26",x"4d",x"26"),
  1890 => (x"4f",x"26",x"4b",x"26"),
  1891 => (x"00",x"00",x"00",x"00"),
  1892 => (x"00",x"00",x"00",x"00"),
  1893 => (x"49",x"4a",x"71",x"1e"),
  1894 => (x"26",x"87",x"eb",x"fc"),
  1895 => (x"4a",x"c0",x"1e",x"4f"),
  1896 => (x"91",x"c4",x"49",x"72"),
  1897 => (x"81",x"ec",x"f7",x"c1"),
  1898 => (x"82",x"c1",x"79",x"c0"),
  1899 => (x"04",x"aa",x"b7",x"d0"),
  1900 => (x"4f",x"26",x"87",x"ee"),
  1901 => (x"5c",x"5b",x"5e",x"0e"),
  1902 => (x"4d",x"71",x"0e",x"5d"),
  1903 => (x"75",x"87",x"cb",x"f8"),
  1904 => (x"2a",x"b7",x"c4",x"4a"),
  1905 => (x"ec",x"f7",x"c1",x"92"),
  1906 => (x"cf",x"4c",x"75",x"82"),
  1907 => (x"6a",x"94",x"c2",x"9c"),
  1908 => (x"2b",x"74",x"4b",x"49"),
  1909 => (x"48",x"c2",x"9b",x"c3"),
  1910 => (x"4c",x"70",x"30",x"74"),
  1911 => (x"48",x"74",x"bc",x"ff"),
  1912 => (x"7a",x"70",x"98",x"71"),
  1913 => (x"73",x"87",x"db",x"f7"),
  1914 => (x"87",x"d8",x"fe",x"48"),
  1915 => (x"00",x"00",x"00",x"00"),
  1916 => (x"00",x"00",x"00",x"00"),
  1917 => (x"00",x"00",x"00",x"00"),
  1918 => (x"00",x"00",x"00",x"00"),
  1919 => (x"00",x"00",x"00",x"00"),
  1920 => (x"00",x"00",x"00",x"00"),
  1921 => (x"00",x"00",x"00",x"00"),
  1922 => (x"00",x"00",x"00",x"00"),
  1923 => (x"00",x"00",x"00",x"00"),
  1924 => (x"00",x"00",x"00",x"00"),
  1925 => (x"00",x"00",x"00",x"00"),
  1926 => (x"00",x"00",x"00",x"00"),
  1927 => (x"00",x"00",x"00",x"00"),
  1928 => (x"00",x"00",x"00",x"00"),
  1929 => (x"00",x"00",x"00",x"00"),
  1930 => (x"00",x"00",x"00",x"00"),
  1931 => (x"48",x"d0",x"ff",x"1e"),
  1932 => (x"71",x"78",x"e1",x"c8"),
  1933 => (x"08",x"d4",x"ff",x"48"),
  1934 => (x"48",x"66",x"c4",x"78"),
  1935 => (x"78",x"08",x"d4",x"ff"),
  1936 => (x"71",x"1e",x"4f",x"26"),
  1937 => (x"49",x"66",x"c4",x"4a"),
  1938 => (x"ff",x"49",x"72",x"1e"),
  1939 => (x"d0",x"ff",x"87",x"de"),
  1940 => (x"78",x"e0",x"c0",x"48"),
  1941 => (x"1e",x"4f",x"26",x"26"),
  1942 => (x"4b",x"71",x"1e",x"73"),
  1943 => (x"1e",x"49",x"66",x"c8"),
  1944 => (x"e0",x"c1",x"4a",x"73"),
  1945 => (x"d9",x"ff",x"49",x"a2"),
  1946 => (x"87",x"c4",x"26",x"87"),
  1947 => (x"4c",x"26",x"4d",x"26"),
  1948 => (x"4f",x"26",x"4b",x"26"),
  1949 => (x"4a",x"d4",x"ff",x"1e"),
  1950 => (x"ff",x"7a",x"ff",x"c3"),
  1951 => (x"e1",x"c8",x"48",x"d0"),
  1952 => (x"c3",x"7a",x"de",x"78"),
  1953 => (x"7a",x"bf",x"c8",x"e3"),
  1954 => (x"28",x"c8",x"48",x"49"),
  1955 => (x"48",x"71",x"7a",x"70"),
  1956 => (x"7a",x"70",x"28",x"d0"),
  1957 => (x"28",x"d8",x"48",x"71"),
  1958 => (x"d0",x"ff",x"7a",x"70"),
  1959 => (x"78",x"e0",x"c0",x"48"),
  1960 => (x"5e",x"0e",x"4f",x"26"),
  1961 => (x"0e",x"5d",x"5c",x"5b"),
  1962 => (x"e3",x"c3",x"4c",x"71"),
  1963 => (x"4b",x"4d",x"bf",x"c8"),
  1964 => (x"66",x"d0",x"2b",x"74"),
  1965 => (x"d4",x"83",x"c1",x"9b"),
  1966 => (x"c2",x"04",x"ab",x"66"),
  1967 => (x"74",x"4b",x"c0",x"87"),
  1968 => (x"49",x"66",x"d0",x"4a"),
  1969 => (x"b9",x"ff",x"31",x"72"),
  1970 => (x"48",x"73",x"99",x"75"),
  1971 => (x"4a",x"70",x"30",x"72"),
  1972 => (x"c3",x"b0",x"71",x"48"),
  1973 => (x"fe",x"58",x"cc",x"e3"),
  1974 => (x"4d",x"26",x"87",x"da"),
  1975 => (x"4b",x"26",x"4c",x"26"),
  1976 => (x"5e",x"0e",x"4f",x"26"),
  1977 => (x"0e",x"5d",x"5c",x"5b"),
  1978 => (x"c3",x"4c",x"71",x"1e"),
  1979 => (x"c0",x"4b",x"cc",x"e3"),
  1980 => (x"49",x"f4",x"c0",x"4a"),
  1981 => (x"87",x"cd",x"c7",x"fe"),
  1982 => (x"e3",x"c3",x"1e",x"74"),
  1983 => (x"e7",x"fe",x"49",x"cc"),
  1984 => (x"86",x"c4",x"87",x"df"),
  1985 => (x"02",x"99",x"49",x"70"),
  1986 => (x"c4",x"87",x"ea",x"c0"),
  1987 => (x"1e",x"4d",x"a6",x"1e"),
  1988 => (x"49",x"cc",x"e3",x"c3"),
  1989 => (x"87",x"e3",x"ee",x"fe"),
  1990 => (x"98",x"70",x"86",x"c8"),
  1991 => (x"75",x"87",x"d6",x"02"),
  1992 => (x"eb",x"fd",x"c1",x"4a"),
  1993 => (x"fe",x"4b",x"c4",x"49"),
  1994 => (x"70",x"87",x"ff",x"c4"),
  1995 => (x"87",x"ca",x"02",x"98"),
  1996 => (x"ed",x"c0",x"48",x"c0"),
  1997 => (x"c0",x"48",x"c0",x"87"),
  1998 => (x"f3",x"c0",x"87",x"e8"),
  1999 => (x"87",x"c4",x"c1",x"87"),
  2000 => (x"c8",x"02",x"98",x"70"),
  2001 => (x"87",x"fc",x"c0",x"87"),
  2002 => (x"f8",x"05",x"98",x"70"),
  2003 => (x"ec",x"e3",x"c3",x"87"),
  2004 => (x"87",x"cc",x"02",x"bf"),
  2005 => (x"48",x"c8",x"e3",x"c3"),
  2006 => (x"bf",x"ec",x"e3",x"c3"),
  2007 => (x"87",x"d4",x"fc",x"78"),
  2008 => (x"26",x"26",x"48",x"c1"),
  2009 => (x"26",x"4c",x"26",x"4d"),
  2010 => (x"5b",x"4f",x"26",x"4b"),
  2011 => (x"00",x"43",x"52",x"41"),
  2012 => (x"c3",x"1e",x"c0",x"1e"),
  2013 => (x"fe",x"49",x"cc",x"e3"),
  2014 => (x"c3",x"87",x"d9",x"eb"),
  2015 => (x"c0",x"48",x"e4",x"e3"),
  2016 => (x"4f",x"26",x"26",x"78"),
  2017 => (x"5c",x"5b",x"5e",x"0e"),
  2018 => (x"86",x"f4",x"0e",x"5d"),
  2019 => (x"c0",x"48",x"a6",x"c4"),
  2020 => (x"e4",x"e3",x"c3",x"78"),
  2021 => (x"b7",x"c3",x"48",x"bf"),
  2022 => (x"87",x"d1",x"03",x"a8"),
  2023 => (x"bf",x"e4",x"e3",x"c3"),
  2024 => (x"c3",x"80",x"c1",x"48"),
  2025 => (x"c0",x"58",x"e8",x"e3"),
  2026 => (x"e2",x"c6",x"48",x"fb"),
  2027 => (x"cc",x"e3",x"c3",x"87"),
  2028 => (x"da",x"f0",x"fe",x"49"),
  2029 => (x"c3",x"4c",x"70",x"87"),
  2030 => (x"4a",x"bf",x"e4",x"e3"),
  2031 => (x"d8",x"02",x"8a",x"c3"),
  2032 => (x"02",x"8a",x"c1",x"87"),
  2033 => (x"8a",x"87",x"cb",x"c5"),
  2034 => (x"87",x"f6",x"c2",x"02"),
  2035 => (x"cd",x"c1",x"02",x"8a"),
  2036 => (x"c3",x"02",x"8a",x"87"),
  2037 => (x"e1",x"c5",x"87",x"e2"),
  2038 => (x"75",x"4d",x"c0",x"87"),
  2039 => (x"c2",x"92",x"c4",x"4a"),
  2040 => (x"c3",x"82",x"ed",x"c5"),
  2041 => (x"75",x"48",x"e0",x"e3"),
  2042 => (x"6e",x"7e",x"70",x"80"),
  2043 => (x"49",x"4b",x"bf",x"97"),
  2044 => (x"c1",x"48",x"6e",x"4b"),
  2045 => (x"81",x"6a",x"50",x"a3"),
  2046 => (x"a6",x"cc",x"48",x"11"),
  2047 => (x"02",x"ac",x"70",x"58"),
  2048 => (x"48",x"6e",x"87",x"c4"),
  2049 => (x"66",x"c8",x"50",x"c0"),
  2050 => (x"c3",x"87",x"c7",x"05"),
  2051 => (x"c4",x"48",x"e4",x"e3"),
  2052 => (x"85",x"c1",x"78",x"a5"),
  2053 => (x"04",x"ad",x"b7",x"c4"),
  2054 => (x"c4",x"87",x"c0",x"ff"),
  2055 => (x"e3",x"c3",x"87",x"dc"),
  2056 => (x"c8",x"48",x"bf",x"f0"),
  2057 => (x"d1",x"01",x"a8",x"b7"),
  2058 => (x"02",x"ac",x"ca",x"87"),
  2059 => (x"ac",x"cd",x"87",x"cc"),
  2060 => (x"c0",x"87",x"c7",x"02"),
  2061 => (x"c0",x"03",x"ac",x"b7"),
  2062 => (x"e3",x"c3",x"87",x"f3"),
  2063 => (x"c8",x"4b",x"bf",x"f0"),
  2064 => (x"d2",x"03",x"ab",x"b7"),
  2065 => (x"f4",x"e3",x"c3",x"87"),
  2066 => (x"c0",x"81",x"73",x"49"),
  2067 => (x"83",x"c1",x"51",x"e0"),
  2068 => (x"04",x"ab",x"b7",x"c8"),
  2069 => (x"c3",x"87",x"ee",x"ff"),
  2070 => (x"c1",x"48",x"fc",x"e3"),
  2071 => (x"cf",x"c1",x"50",x"d2"),
  2072 => (x"50",x"cd",x"c1",x"50"),
  2073 => (x"80",x"e4",x"50",x"c0"),
  2074 => (x"cd",x"c3",x"78",x"c3"),
  2075 => (x"f0",x"e3",x"c3",x"87"),
  2076 => (x"c1",x"48",x"49",x"bf"),
  2077 => (x"f4",x"e3",x"c3",x"80"),
  2078 => (x"a0",x"c4",x"48",x"58"),
  2079 => (x"c2",x"51",x"74",x"81"),
  2080 => (x"f0",x"c0",x"87",x"f8"),
  2081 => (x"da",x"04",x"ac",x"b7"),
  2082 => (x"b7",x"f9",x"c0",x"87"),
  2083 => (x"87",x"d3",x"01",x"ac"),
  2084 => (x"bf",x"e8",x"e3",x"c3"),
  2085 => (x"74",x"91",x"ca",x"49"),
  2086 => (x"8a",x"f0",x"c0",x"4a"),
  2087 => (x"48",x"e8",x"e3",x"c3"),
  2088 => (x"ca",x"78",x"a1",x"72"),
  2089 => (x"c6",x"c0",x"02",x"ac"),
  2090 => (x"05",x"ac",x"cd",x"87"),
  2091 => (x"c3",x"87",x"cb",x"c2"),
  2092 => (x"c3",x"48",x"e4",x"e3"),
  2093 => (x"87",x"c2",x"c2",x"78"),
  2094 => (x"ac",x"b7",x"f0",x"c0"),
  2095 => (x"c0",x"87",x"db",x"04"),
  2096 => (x"01",x"ac",x"b7",x"f9"),
  2097 => (x"c3",x"87",x"d3",x"c0"),
  2098 => (x"49",x"bf",x"ec",x"e3"),
  2099 => (x"4a",x"74",x"91",x"d0"),
  2100 => (x"c3",x"8a",x"f0",x"c0"),
  2101 => (x"72",x"48",x"ec",x"e3"),
  2102 => (x"c1",x"c1",x"78",x"a1"),
  2103 => (x"c0",x"04",x"ac",x"b7"),
  2104 => (x"c6",x"c1",x"87",x"db"),
  2105 => (x"c0",x"01",x"ac",x"b7"),
  2106 => (x"e3",x"c3",x"87",x"d3"),
  2107 => (x"d0",x"49",x"bf",x"ec"),
  2108 => (x"c0",x"4a",x"74",x"91"),
  2109 => (x"e3",x"c3",x"8a",x"f7"),
  2110 => (x"a1",x"72",x"48",x"ec"),
  2111 => (x"02",x"ac",x"ca",x"78"),
  2112 => (x"cd",x"87",x"c6",x"c0"),
  2113 => (x"f1",x"c0",x"05",x"ac"),
  2114 => (x"e4",x"e3",x"c3",x"87"),
  2115 => (x"c0",x"78",x"c3",x"48"),
  2116 => (x"e2",x"c0",x"87",x"e8"),
  2117 => (x"c9",x"c0",x"05",x"ac"),
  2118 => (x"48",x"a6",x"c4",x"87"),
  2119 => (x"c0",x"78",x"fb",x"c0"),
  2120 => (x"ac",x"ca",x"87",x"d8"),
  2121 => (x"87",x"c6",x"c0",x"02"),
  2122 => (x"c0",x"05",x"ac",x"cd"),
  2123 => (x"e3",x"c3",x"87",x"c9"),
  2124 => (x"78",x"c3",x"48",x"e4"),
  2125 => (x"c8",x"87",x"c3",x"c0"),
  2126 => (x"b7",x"c0",x"5c",x"a6"),
  2127 => (x"c4",x"c0",x"03",x"ac"),
  2128 => (x"ca",x"c0",x"48",x"87"),
  2129 => (x"02",x"66",x"c4",x"87"),
  2130 => (x"48",x"87",x"c6",x"f9"),
  2131 => (x"f4",x"99",x"ff",x"c3"),
  2132 => (x"87",x"cf",x"f8",x"8e"),
  2133 => (x"46",x"4e",x"4f",x"43"),
  2134 => (x"4f",x"4d",x"00",x"3d"),
  2135 => (x"41",x"4e",x"00",x"44"),
  2136 => (x"44",x"00",x"45",x"4d"),
  2137 => (x"55",x"41",x"46",x"45"),
  2138 => (x"30",x"3d",x"54",x"4c"),
  2139 => (x"00",x"21",x"54",x"00"),
  2140 => (x"00",x"21",x"5a",x"00"),
  2141 => (x"00",x"21",x"5e",x"00"),
  2142 => (x"00",x"21",x"63",x"00"),
  2143 => (x"d0",x"ff",x"1e",x"00"),
  2144 => (x"78",x"c9",x"c8",x"48"),
  2145 => (x"d4",x"ff",x"48",x"71"),
  2146 => (x"4f",x"26",x"78",x"08"),
  2147 => (x"49",x"4a",x"71",x"1e"),
  2148 => (x"d0",x"ff",x"87",x"eb"),
  2149 => (x"26",x"78",x"c8",x"48"),
  2150 => (x"1e",x"73",x"1e",x"4f"),
  2151 => (x"e4",x"c3",x"4b",x"71"),
  2152 => (x"c3",x"02",x"bf",x"cc"),
  2153 => (x"87",x"eb",x"c2",x"87"),
  2154 => (x"c8",x"48",x"d0",x"ff"),
  2155 => (x"49",x"73",x"78",x"c9"),
  2156 => (x"ff",x"b1",x"e0",x"c0"),
  2157 => (x"78",x"71",x"48",x"d4"),
  2158 => (x"48",x"c0",x"e4",x"c3"),
  2159 => (x"66",x"c8",x"78",x"c0"),
  2160 => (x"c3",x"87",x"c5",x"02"),
  2161 => (x"87",x"c2",x"49",x"ff"),
  2162 => (x"e4",x"c3",x"49",x"c0"),
  2163 => (x"66",x"cc",x"59",x"c8"),
  2164 => (x"c5",x"87",x"c6",x"02"),
  2165 => (x"c4",x"4a",x"d5",x"d5"),
  2166 => (x"ff",x"ff",x"cf",x"87"),
  2167 => (x"cc",x"e4",x"c3",x"4a"),
  2168 => (x"cc",x"e4",x"c3",x"5a"),
  2169 => (x"c4",x"78",x"c1",x"48"),
  2170 => (x"26",x"4d",x"26",x"87"),
  2171 => (x"26",x"4b",x"26",x"4c"),
  2172 => (x"5b",x"5e",x"0e",x"4f"),
  2173 => (x"71",x"0e",x"5d",x"5c"),
  2174 => (x"c8",x"e4",x"c3",x"4a"),
  2175 => (x"9a",x"72",x"4c",x"bf"),
  2176 => (x"49",x"87",x"cb",x"02"),
  2177 => (x"c6",x"c2",x"91",x"c8"),
  2178 => (x"83",x"71",x"4b",x"cf"),
  2179 => (x"ca",x"c2",x"87",x"c4"),
  2180 => (x"4d",x"c0",x"4b",x"cf"),
  2181 => (x"99",x"74",x"49",x"13"),
  2182 => (x"bf",x"c4",x"e4",x"c3"),
  2183 => (x"48",x"d4",x"ff",x"b9"),
  2184 => (x"b7",x"c1",x"78",x"71"),
  2185 => (x"b7",x"c8",x"85",x"2c"),
  2186 => (x"87",x"e8",x"04",x"ad"),
  2187 => (x"bf",x"c0",x"e4",x"c3"),
  2188 => (x"c3",x"80",x"c8",x"48"),
  2189 => (x"fe",x"58",x"c4",x"e4"),
  2190 => (x"73",x"1e",x"87",x"ef"),
  2191 => (x"13",x"4b",x"71",x"1e"),
  2192 => (x"cb",x"02",x"9a",x"4a"),
  2193 => (x"fe",x"49",x"72",x"87"),
  2194 => (x"4a",x"13",x"87",x"e7"),
  2195 => (x"87",x"f5",x"05",x"9a"),
  2196 => (x"1e",x"87",x"da",x"fe"),
  2197 => (x"bf",x"c0",x"e4",x"c3"),
  2198 => (x"c0",x"e4",x"c3",x"49"),
  2199 => (x"78",x"a1",x"c1",x"48"),
  2200 => (x"a9",x"b7",x"c0",x"c4"),
  2201 => (x"ff",x"87",x"db",x"03"),
  2202 => (x"e4",x"c3",x"48",x"d4"),
  2203 => (x"c3",x"78",x"bf",x"c4"),
  2204 => (x"49",x"bf",x"c0",x"e4"),
  2205 => (x"48",x"c0",x"e4",x"c3"),
  2206 => (x"c4",x"78",x"a1",x"c1"),
  2207 => (x"04",x"a9",x"b7",x"c0"),
  2208 => (x"d0",x"ff",x"87",x"e5"),
  2209 => (x"c3",x"78",x"c8",x"48"),
  2210 => (x"c0",x"48",x"cc",x"e4"),
  2211 => (x"00",x"4f",x"26",x"78"),
  2212 => (x"00",x"00",x"00",x"00"),
  2213 => (x"00",x"00",x"00",x"00"),
  2214 => (x"5f",x"5f",x"00",x"00"),
  2215 => (x"00",x"00",x"00",x"00"),
  2216 => (x"03",x"00",x"03",x"03"),
  2217 => (x"14",x"00",x"00",x"03"),
  2218 => (x"7f",x"14",x"7f",x"7f"),
  2219 => (x"00",x"00",x"14",x"7f"),
  2220 => (x"6b",x"6b",x"2e",x"24"),
  2221 => (x"4c",x"00",x"12",x"3a"),
  2222 => (x"6c",x"18",x"36",x"6a"),
  2223 => (x"30",x"00",x"32",x"56"),
  2224 => (x"77",x"59",x"4f",x"7e"),
  2225 => (x"00",x"40",x"68",x"3a"),
  2226 => (x"03",x"07",x"04",x"00"),
  2227 => (x"00",x"00",x"00",x"00"),
  2228 => (x"63",x"3e",x"1c",x"00"),
  2229 => (x"00",x"00",x"00",x"41"),
  2230 => (x"3e",x"63",x"41",x"00"),
  2231 => (x"08",x"00",x"00",x"1c"),
  2232 => (x"1c",x"1c",x"3e",x"2a"),
  2233 => (x"00",x"08",x"2a",x"3e"),
  2234 => (x"3e",x"3e",x"08",x"08"),
  2235 => (x"00",x"00",x"08",x"08"),
  2236 => (x"60",x"e0",x"80",x"00"),
  2237 => (x"00",x"00",x"00",x"00"),
  2238 => (x"08",x"08",x"08",x"08"),
  2239 => (x"00",x"00",x"08",x"08"),
  2240 => (x"60",x"60",x"00",x"00"),
  2241 => (x"40",x"00",x"00",x"00"),
  2242 => (x"0c",x"18",x"30",x"60"),
  2243 => (x"00",x"01",x"03",x"06"),
  2244 => (x"4d",x"59",x"7f",x"3e"),
  2245 => (x"00",x"00",x"3e",x"7f"),
  2246 => (x"7f",x"7f",x"06",x"04"),
  2247 => (x"00",x"00",x"00",x"00"),
  2248 => (x"59",x"71",x"63",x"42"),
  2249 => (x"00",x"00",x"46",x"4f"),
  2250 => (x"49",x"49",x"63",x"22"),
  2251 => (x"18",x"00",x"36",x"7f"),
  2252 => (x"7f",x"13",x"16",x"1c"),
  2253 => (x"00",x"00",x"10",x"7f"),
  2254 => (x"45",x"45",x"67",x"27"),
  2255 => (x"00",x"00",x"39",x"7d"),
  2256 => (x"49",x"4b",x"7e",x"3c"),
  2257 => (x"00",x"00",x"30",x"79"),
  2258 => (x"79",x"71",x"01",x"01"),
  2259 => (x"00",x"00",x"07",x"0f"),
  2260 => (x"49",x"49",x"7f",x"36"),
  2261 => (x"00",x"00",x"36",x"7f"),
  2262 => (x"69",x"49",x"4f",x"06"),
  2263 => (x"00",x"00",x"1e",x"3f"),
  2264 => (x"66",x"66",x"00",x"00"),
  2265 => (x"00",x"00",x"00",x"00"),
  2266 => (x"66",x"e6",x"80",x"00"),
  2267 => (x"00",x"00",x"00",x"00"),
  2268 => (x"14",x"14",x"08",x"08"),
  2269 => (x"00",x"00",x"22",x"22"),
  2270 => (x"14",x"14",x"14",x"14"),
  2271 => (x"00",x"00",x"14",x"14"),
  2272 => (x"14",x"14",x"22",x"22"),
  2273 => (x"00",x"00",x"08",x"08"),
  2274 => (x"59",x"51",x"03",x"02"),
  2275 => (x"3e",x"00",x"06",x"0f"),
  2276 => (x"55",x"5d",x"41",x"7f"),
  2277 => (x"00",x"00",x"1e",x"1f"),
  2278 => (x"09",x"09",x"7f",x"7e"),
  2279 => (x"00",x"00",x"7e",x"7f"),
  2280 => (x"49",x"49",x"7f",x"7f"),
  2281 => (x"00",x"00",x"36",x"7f"),
  2282 => (x"41",x"63",x"3e",x"1c"),
  2283 => (x"00",x"00",x"41",x"41"),
  2284 => (x"63",x"41",x"7f",x"7f"),
  2285 => (x"00",x"00",x"1c",x"3e"),
  2286 => (x"49",x"49",x"7f",x"7f"),
  2287 => (x"00",x"00",x"41",x"41"),
  2288 => (x"09",x"09",x"7f",x"7f"),
  2289 => (x"00",x"00",x"01",x"01"),
  2290 => (x"49",x"41",x"7f",x"3e"),
  2291 => (x"00",x"00",x"7a",x"7b"),
  2292 => (x"08",x"08",x"7f",x"7f"),
  2293 => (x"00",x"00",x"7f",x"7f"),
  2294 => (x"7f",x"7f",x"41",x"00"),
  2295 => (x"00",x"00",x"00",x"41"),
  2296 => (x"40",x"40",x"60",x"20"),
  2297 => (x"7f",x"00",x"3f",x"7f"),
  2298 => (x"36",x"1c",x"08",x"7f"),
  2299 => (x"00",x"00",x"41",x"63"),
  2300 => (x"40",x"40",x"7f",x"7f"),
  2301 => (x"7f",x"00",x"40",x"40"),
  2302 => (x"06",x"0c",x"06",x"7f"),
  2303 => (x"7f",x"00",x"7f",x"7f"),
  2304 => (x"18",x"0c",x"06",x"7f"),
  2305 => (x"00",x"00",x"7f",x"7f"),
  2306 => (x"41",x"41",x"7f",x"3e"),
  2307 => (x"00",x"00",x"3e",x"7f"),
  2308 => (x"09",x"09",x"7f",x"7f"),
  2309 => (x"3e",x"00",x"06",x"0f"),
  2310 => (x"7f",x"61",x"41",x"7f"),
  2311 => (x"00",x"00",x"40",x"7e"),
  2312 => (x"19",x"09",x"7f",x"7f"),
  2313 => (x"00",x"00",x"66",x"7f"),
  2314 => (x"59",x"4d",x"6f",x"26"),
  2315 => (x"00",x"00",x"32",x"7b"),
  2316 => (x"7f",x"7f",x"01",x"01"),
  2317 => (x"00",x"00",x"01",x"01"),
  2318 => (x"40",x"40",x"7f",x"3f"),
  2319 => (x"00",x"00",x"3f",x"7f"),
  2320 => (x"70",x"70",x"3f",x"0f"),
  2321 => (x"7f",x"00",x"0f",x"3f"),
  2322 => (x"30",x"18",x"30",x"7f"),
  2323 => (x"41",x"00",x"7f",x"7f"),
  2324 => (x"1c",x"1c",x"36",x"63"),
  2325 => (x"01",x"41",x"63",x"36"),
  2326 => (x"7c",x"7c",x"06",x"03"),
  2327 => (x"61",x"01",x"03",x"06"),
  2328 => (x"47",x"4d",x"59",x"71"),
  2329 => (x"00",x"00",x"41",x"43"),
  2330 => (x"41",x"7f",x"7f",x"00"),
  2331 => (x"01",x"00",x"00",x"41"),
  2332 => (x"18",x"0c",x"06",x"03"),
  2333 => (x"00",x"40",x"60",x"30"),
  2334 => (x"7f",x"41",x"41",x"00"),
  2335 => (x"08",x"00",x"00",x"7f"),
  2336 => (x"06",x"03",x"06",x"0c"),
  2337 => (x"80",x"00",x"08",x"0c"),
  2338 => (x"80",x"80",x"80",x"80"),
  2339 => (x"00",x"00",x"80",x"80"),
  2340 => (x"07",x"03",x"00",x"00"),
  2341 => (x"00",x"00",x"00",x"04"),
  2342 => (x"54",x"54",x"74",x"20"),
  2343 => (x"00",x"00",x"78",x"7c"),
  2344 => (x"44",x"44",x"7f",x"7f"),
  2345 => (x"00",x"00",x"38",x"7c"),
  2346 => (x"44",x"44",x"7c",x"38"),
  2347 => (x"00",x"00",x"00",x"44"),
  2348 => (x"44",x"44",x"7c",x"38"),
  2349 => (x"00",x"00",x"7f",x"7f"),
  2350 => (x"54",x"54",x"7c",x"38"),
  2351 => (x"00",x"00",x"18",x"5c"),
  2352 => (x"05",x"7f",x"7e",x"04"),
  2353 => (x"00",x"00",x"00",x"05"),
  2354 => (x"a4",x"a4",x"bc",x"18"),
  2355 => (x"00",x"00",x"7c",x"fc"),
  2356 => (x"04",x"04",x"7f",x"7f"),
  2357 => (x"00",x"00",x"78",x"7c"),
  2358 => (x"7d",x"3d",x"00",x"00"),
  2359 => (x"00",x"00",x"00",x"40"),
  2360 => (x"fd",x"80",x"80",x"80"),
  2361 => (x"00",x"00",x"00",x"7d"),
  2362 => (x"38",x"10",x"7f",x"7f"),
  2363 => (x"00",x"00",x"44",x"6c"),
  2364 => (x"7f",x"3f",x"00",x"00"),
  2365 => (x"7c",x"00",x"00",x"40"),
  2366 => (x"0c",x"18",x"0c",x"7c"),
  2367 => (x"00",x"00",x"78",x"7c"),
  2368 => (x"04",x"04",x"7c",x"7c"),
  2369 => (x"00",x"00",x"78",x"7c"),
  2370 => (x"44",x"44",x"7c",x"38"),
  2371 => (x"00",x"00",x"38",x"7c"),
  2372 => (x"24",x"24",x"fc",x"fc"),
  2373 => (x"00",x"00",x"18",x"3c"),
  2374 => (x"24",x"24",x"3c",x"18"),
  2375 => (x"00",x"00",x"fc",x"fc"),
  2376 => (x"04",x"04",x"7c",x"7c"),
  2377 => (x"00",x"00",x"08",x"0c"),
  2378 => (x"54",x"54",x"5c",x"48"),
  2379 => (x"00",x"00",x"20",x"74"),
  2380 => (x"44",x"7f",x"3f",x"04"),
  2381 => (x"00",x"00",x"00",x"44"),
  2382 => (x"40",x"40",x"7c",x"3c"),
  2383 => (x"00",x"00",x"7c",x"7c"),
  2384 => (x"60",x"60",x"3c",x"1c"),
  2385 => (x"3c",x"00",x"1c",x"3c"),
  2386 => (x"60",x"30",x"60",x"7c"),
  2387 => (x"44",x"00",x"3c",x"7c"),
  2388 => (x"38",x"10",x"38",x"6c"),
  2389 => (x"00",x"00",x"44",x"6c"),
  2390 => (x"60",x"e0",x"bc",x"1c"),
  2391 => (x"00",x"00",x"1c",x"3c"),
  2392 => (x"5c",x"74",x"64",x"44"),
  2393 => (x"00",x"00",x"44",x"4c"),
  2394 => (x"77",x"3e",x"08",x"08"),
  2395 => (x"00",x"00",x"41",x"41"),
  2396 => (x"7f",x"7f",x"00",x"00"),
  2397 => (x"00",x"00",x"00",x"00"),
  2398 => (x"3e",x"77",x"41",x"41"),
  2399 => (x"02",x"00",x"08",x"08"),
  2400 => (x"02",x"03",x"01",x"01"),
  2401 => (x"7f",x"00",x"01",x"02"),
  2402 => (x"7f",x"7f",x"7f",x"7f"),
  2403 => (x"08",x"00",x"7f",x"7f"),
  2404 => (x"3e",x"1c",x"1c",x"08"),
  2405 => (x"7f",x"7f",x"7f",x"3e"),
  2406 => (x"1c",x"3e",x"3e",x"7f"),
  2407 => (x"00",x"08",x"08",x"1c"),
  2408 => (x"7c",x"7c",x"18",x"10"),
  2409 => (x"00",x"00",x"10",x"18"),
  2410 => (x"7c",x"7c",x"30",x"10"),
  2411 => (x"10",x"00",x"10",x"30"),
  2412 => (x"78",x"60",x"60",x"30"),
  2413 => (x"42",x"00",x"06",x"1e"),
  2414 => (x"3c",x"18",x"3c",x"66"),
  2415 => (x"78",x"00",x"42",x"66"),
  2416 => (x"c6",x"c2",x"6a",x"38"),
  2417 => (x"60",x"00",x"38",x"6c"),
  2418 => (x"00",x"60",x"00",x"00"),
  2419 => (x"0e",x"00",x"60",x"00"),
  2420 => (x"5d",x"5c",x"5b",x"5e"),
  2421 => (x"4c",x"71",x"1e",x"0e"),
  2422 => (x"bf",x"dd",x"e4",x"c3"),
  2423 => (x"c0",x"4b",x"c0",x"4d"),
  2424 => (x"02",x"ab",x"74",x"1e"),
  2425 => (x"a6",x"c4",x"87",x"c7"),
  2426 => (x"c5",x"78",x"c0",x"48"),
  2427 => (x"48",x"a6",x"c4",x"87"),
  2428 => (x"66",x"c4",x"78",x"c1"),
  2429 => (x"ee",x"49",x"73",x"1e"),
  2430 => (x"86",x"c8",x"87",x"df"),
  2431 => (x"ef",x"49",x"e0",x"c0"),
  2432 => (x"a5",x"c4",x"87",x"ef"),
  2433 => (x"f0",x"49",x"6a",x"4a"),
  2434 => (x"c6",x"f1",x"87",x"f0"),
  2435 => (x"c1",x"85",x"cb",x"87"),
  2436 => (x"ab",x"b7",x"c8",x"83"),
  2437 => (x"87",x"c7",x"ff",x"04"),
  2438 => (x"26",x"4d",x"26",x"26"),
  2439 => (x"26",x"4b",x"26",x"4c"),
  2440 => (x"4a",x"71",x"1e",x"4f"),
  2441 => (x"5a",x"e1",x"e4",x"c3"),
  2442 => (x"48",x"e1",x"e4",x"c3"),
  2443 => (x"fe",x"49",x"78",x"c7"),
  2444 => (x"4f",x"26",x"87",x"dd"),
  2445 => (x"71",x"1e",x"73",x"1e"),
  2446 => (x"aa",x"b7",x"c0",x"4a"),
  2447 => (x"c2",x"87",x"d3",x"03"),
  2448 => (x"05",x"bf",x"d7",x"e6"),
  2449 => (x"4b",x"c1",x"87",x"c4"),
  2450 => (x"4b",x"c0",x"87",x"c2"),
  2451 => (x"5b",x"db",x"e6",x"c2"),
  2452 => (x"e6",x"c2",x"87",x"c4"),
  2453 => (x"e6",x"c2",x"5a",x"db"),
  2454 => (x"c1",x"4a",x"bf",x"d7"),
  2455 => (x"a2",x"c0",x"c1",x"9a"),
  2456 => (x"87",x"e8",x"ec",x"49"),
  2457 => (x"e6",x"c2",x"48",x"fc"),
  2458 => (x"fe",x"78",x"bf",x"d7"),
  2459 => (x"71",x"1e",x"87",x"ef"),
  2460 => (x"1e",x"66",x"c4",x"4a"),
  2461 => (x"df",x"ff",x"49",x"72"),
  2462 => (x"26",x"26",x"87",x"dd"),
  2463 => (x"e6",x"c2",x"1e",x"4f"),
  2464 => (x"ff",x"49",x"bf",x"d7"),
  2465 => (x"c3",x"87",x"cd",x"dc"),
  2466 => (x"e8",x"48",x"d5",x"e4"),
  2467 => (x"e4",x"c3",x"78",x"bf"),
  2468 => (x"bf",x"ec",x"48",x"d1"),
  2469 => (x"d5",x"e4",x"c3",x"78"),
  2470 => (x"c3",x"49",x"4a",x"bf"),
  2471 => (x"b7",x"c8",x"99",x"ff"),
  2472 => (x"71",x"48",x"72",x"2a"),
  2473 => (x"dd",x"e4",x"c3",x"b0"),
  2474 => (x"0e",x"4f",x"26",x"58"),
  2475 => (x"5d",x"5c",x"5b",x"5e"),
  2476 => (x"ff",x"4b",x"71",x"0e"),
  2477 => (x"e4",x"c3",x"87",x"c7"),
  2478 => (x"50",x"c0",x"48",x"d0"),
  2479 => (x"db",x"ff",x"49",x"73"),
  2480 => (x"49",x"70",x"87",x"f2"),
  2481 => (x"cb",x"9c",x"c2",x"4c"),
  2482 => (x"d2",x"cb",x"49",x"ee"),
  2483 => (x"4d",x"49",x"70",x"87"),
  2484 => (x"97",x"d0",x"e4",x"c3"),
  2485 => (x"e4",x"c1",x"05",x"bf"),
  2486 => (x"49",x"66",x"d0",x"87"),
  2487 => (x"bf",x"d9",x"e4",x"c3"),
  2488 => (x"87",x"d7",x"05",x"99"),
  2489 => (x"c3",x"49",x"66",x"d4"),
  2490 => (x"99",x"bf",x"d1",x"e4"),
  2491 => (x"73",x"87",x"cc",x"05"),
  2492 => (x"ff",x"da",x"ff",x"49"),
  2493 => (x"02",x"98",x"70",x"87"),
  2494 => (x"c1",x"87",x"c2",x"c1"),
  2495 => (x"87",x"fd",x"fd",x"4c"),
  2496 => (x"e6",x"ca",x"49",x"75"),
  2497 => (x"02",x"98",x"70",x"87"),
  2498 => (x"e4",x"c3",x"87",x"c6"),
  2499 => (x"50",x"c1",x"48",x"d0"),
  2500 => (x"97",x"d0",x"e4",x"c3"),
  2501 => (x"e4",x"c0",x"05",x"bf"),
  2502 => (x"d9",x"e4",x"c3",x"87"),
  2503 => (x"66",x"d0",x"49",x"bf"),
  2504 => (x"d6",x"ff",x"05",x"99"),
  2505 => (x"d1",x"e4",x"c3",x"87"),
  2506 => (x"66",x"d4",x"49",x"bf"),
  2507 => (x"ca",x"ff",x"05",x"99"),
  2508 => (x"ff",x"49",x"73",x"87"),
  2509 => (x"70",x"87",x"fd",x"d9"),
  2510 => (x"fe",x"fe",x"05",x"98"),
  2511 => (x"fb",x"48",x"74",x"87"),
  2512 => (x"5e",x"0e",x"87",x"d7"),
  2513 => (x"0e",x"5d",x"5c",x"5b"),
  2514 => (x"4d",x"c0",x"86",x"f4"),
  2515 => (x"7e",x"bf",x"ec",x"4c"),
  2516 => (x"c3",x"48",x"a6",x"c4"),
  2517 => (x"78",x"bf",x"dd",x"e4"),
  2518 => (x"1e",x"c0",x"1e",x"c1"),
  2519 => (x"ca",x"fd",x"49",x"c7"),
  2520 => (x"70",x"86",x"c8",x"87"),
  2521 => (x"87",x"ce",x"02",x"98"),
  2522 => (x"c7",x"fb",x"49",x"ff"),
  2523 => (x"49",x"da",x"c1",x"87"),
  2524 => (x"87",x"c0",x"d9",x"ff"),
  2525 => (x"e4",x"c3",x"4d",x"c1"),
  2526 => (x"02",x"bf",x"97",x"d0"),
  2527 => (x"f2",x"c0",x"87",x"c4"),
  2528 => (x"e4",x"c3",x"87",x"d1"),
  2529 => (x"c2",x"4b",x"bf",x"d5"),
  2530 => (x"05",x"bf",x"d7",x"e6"),
  2531 => (x"c3",x"87",x"eb",x"c0"),
  2532 => (x"d8",x"ff",x"49",x"fd"),
  2533 => (x"fa",x"c3",x"87",x"de"),
  2534 => (x"d7",x"d8",x"ff",x"49"),
  2535 => (x"c3",x"49",x"73",x"87"),
  2536 => (x"1e",x"71",x"99",x"ff"),
  2537 => (x"c5",x"fb",x"49",x"c0"),
  2538 => (x"c8",x"49",x"73",x"87"),
  2539 => (x"1e",x"71",x"29",x"b7"),
  2540 => (x"f9",x"fa",x"49",x"c1"),
  2541 => (x"c6",x"86",x"c8",x"87"),
  2542 => (x"e4",x"c3",x"87",x"c3"),
  2543 => (x"9b",x"4b",x"bf",x"d9"),
  2544 => (x"c2",x"87",x"dd",x"02"),
  2545 => (x"49",x"bf",x"d3",x"e6"),
  2546 => (x"70",x"87",x"e0",x"c7"),
  2547 => (x"87",x"c4",x"05",x"98"),
  2548 => (x"87",x"d2",x"4b",x"c0"),
  2549 => (x"c7",x"49",x"e0",x"c2"),
  2550 => (x"e6",x"c2",x"87",x"c5"),
  2551 => (x"87",x"c6",x"58",x"d7"),
  2552 => (x"48",x"d3",x"e6",x"c2"),
  2553 => (x"49",x"73",x"78",x"c0"),
  2554 => (x"ce",x"05",x"99",x"c2"),
  2555 => (x"49",x"eb",x"c3",x"87"),
  2556 => (x"87",x"c0",x"d7",x"ff"),
  2557 => (x"99",x"c2",x"49",x"70"),
  2558 => (x"fb",x"87",x"c2",x"02"),
  2559 => (x"c1",x"49",x"73",x"4c"),
  2560 => (x"87",x"cf",x"05",x"99"),
  2561 => (x"ff",x"49",x"f4",x"c3"),
  2562 => (x"70",x"87",x"e9",x"d6"),
  2563 => (x"02",x"99",x"c2",x"49"),
  2564 => (x"fa",x"87",x"c2",x"c0"),
  2565 => (x"c8",x"49",x"73",x"4c"),
  2566 => (x"87",x"ce",x"05",x"99"),
  2567 => (x"ff",x"49",x"f5",x"c3"),
  2568 => (x"70",x"87",x"d1",x"d6"),
  2569 => (x"02",x"99",x"c2",x"49"),
  2570 => (x"e4",x"c3",x"87",x"d6"),
  2571 => (x"c0",x"02",x"bf",x"e1"),
  2572 => (x"c1",x"48",x"87",x"ca"),
  2573 => (x"e5",x"e4",x"c3",x"88"),
  2574 => (x"87",x"c2",x"c0",x"58"),
  2575 => (x"4d",x"c1",x"4c",x"ff"),
  2576 => (x"99",x"c4",x"49",x"73"),
  2577 => (x"c3",x"87",x"ce",x"05"),
  2578 => (x"d5",x"ff",x"49",x"f2"),
  2579 => (x"49",x"70",x"87",x"e6"),
  2580 => (x"dc",x"02",x"99",x"c2"),
  2581 => (x"e1",x"e4",x"c3",x"87"),
  2582 => (x"c7",x"48",x"7e",x"bf"),
  2583 => (x"c0",x"03",x"a8",x"b7"),
  2584 => (x"48",x"6e",x"87",x"cb"),
  2585 => (x"e4",x"c3",x"80",x"c1"),
  2586 => (x"c2",x"c0",x"58",x"e5"),
  2587 => (x"c1",x"4c",x"fe",x"87"),
  2588 => (x"49",x"fd",x"c3",x"4d"),
  2589 => (x"87",x"fc",x"d4",x"ff"),
  2590 => (x"99",x"c2",x"49",x"70"),
  2591 => (x"87",x"d5",x"c0",x"02"),
  2592 => (x"bf",x"e1",x"e4",x"c3"),
  2593 => (x"87",x"c9",x"c0",x"02"),
  2594 => (x"48",x"e1",x"e4",x"c3"),
  2595 => (x"c2",x"c0",x"78",x"c0"),
  2596 => (x"c1",x"4c",x"fd",x"87"),
  2597 => (x"49",x"fa",x"c3",x"4d"),
  2598 => (x"87",x"d8",x"d4",x"ff"),
  2599 => (x"99",x"c2",x"49",x"70"),
  2600 => (x"87",x"d9",x"c0",x"02"),
  2601 => (x"bf",x"e1",x"e4",x"c3"),
  2602 => (x"a8",x"b7",x"c7",x"48"),
  2603 => (x"87",x"c9",x"c0",x"03"),
  2604 => (x"48",x"e1",x"e4",x"c3"),
  2605 => (x"c2",x"c0",x"78",x"c7"),
  2606 => (x"c1",x"4c",x"fc",x"87"),
  2607 => (x"ac",x"b7",x"c0",x"4d"),
  2608 => (x"87",x"d1",x"c0",x"03"),
  2609 => (x"c1",x"4a",x"66",x"c4"),
  2610 => (x"02",x"6a",x"82",x"d8"),
  2611 => (x"6a",x"87",x"c6",x"c0"),
  2612 => (x"73",x"49",x"74",x"4b"),
  2613 => (x"c3",x"1e",x"c0",x"0f"),
  2614 => (x"da",x"c1",x"1e",x"f0"),
  2615 => (x"87",x"cb",x"f7",x"49"),
  2616 => (x"98",x"70",x"86",x"c8"),
  2617 => (x"87",x"e2",x"c0",x"02"),
  2618 => (x"c3",x"48",x"a6",x"c8"),
  2619 => (x"78",x"bf",x"e1",x"e4"),
  2620 => (x"cb",x"49",x"66",x"c8"),
  2621 => (x"48",x"66",x"c4",x"91"),
  2622 => (x"7e",x"70",x"80",x"71"),
  2623 => (x"c0",x"02",x"bf",x"6e"),
  2624 => (x"bf",x"6e",x"87",x"c8"),
  2625 => (x"49",x"66",x"c8",x"4b"),
  2626 => (x"9d",x"75",x"0f",x"73"),
  2627 => (x"87",x"c8",x"c0",x"02"),
  2628 => (x"bf",x"e1",x"e4",x"c3"),
  2629 => (x"87",x"f7",x"f2",x"49"),
  2630 => (x"bf",x"db",x"e6",x"c2"),
  2631 => (x"87",x"dd",x"c0",x"02"),
  2632 => (x"87",x"c7",x"c2",x"49"),
  2633 => (x"c0",x"02",x"98",x"70"),
  2634 => (x"e4",x"c3",x"87",x"d3"),
  2635 => (x"f2",x"49",x"bf",x"e1"),
  2636 => (x"49",x"c0",x"87",x"dd"),
  2637 => (x"c2",x"87",x"fd",x"f3"),
  2638 => (x"c0",x"48",x"db",x"e6"),
  2639 => (x"f3",x"8e",x"f4",x"78"),
  2640 => (x"5e",x"0e",x"87",x"d7"),
  2641 => (x"0e",x"5d",x"5c",x"5b"),
  2642 => (x"c3",x"4c",x"71",x"1e"),
  2643 => (x"49",x"bf",x"dd",x"e4"),
  2644 => (x"4d",x"a1",x"cd",x"c1"),
  2645 => (x"69",x"81",x"d1",x"c1"),
  2646 => (x"02",x"9c",x"74",x"7e"),
  2647 => (x"a5",x"c4",x"87",x"cf"),
  2648 => (x"c3",x"7b",x"74",x"4b"),
  2649 => (x"49",x"bf",x"dd",x"e4"),
  2650 => (x"6e",x"87",x"f6",x"f2"),
  2651 => (x"05",x"9c",x"74",x"7b"),
  2652 => (x"4b",x"c0",x"87",x"c4"),
  2653 => (x"4b",x"c1",x"87",x"c2"),
  2654 => (x"f7",x"f2",x"49",x"73"),
  2655 => (x"02",x"66",x"d4",x"87"),
  2656 => (x"da",x"49",x"87",x"c7"),
  2657 => (x"c2",x"4a",x"70",x"87"),
  2658 => (x"c2",x"4a",x"c0",x"87"),
  2659 => (x"26",x"5a",x"df",x"e6"),
  2660 => (x"00",x"87",x"c6",x"f2"),
  2661 => (x"00",x"00",x"00",x"00"),
  2662 => (x"00",x"00",x"00",x"00"),
  2663 => (x"1e",x"00",x"00",x"00"),
  2664 => (x"c8",x"ff",x"4a",x"71"),
  2665 => (x"a1",x"72",x"49",x"bf"),
  2666 => (x"1e",x"4f",x"26",x"48"),
  2667 => (x"89",x"bf",x"c8",x"ff"),
  2668 => (x"c0",x"c0",x"c0",x"fe"),
  2669 => (x"01",x"a9",x"c0",x"c0"),
  2670 => (x"4a",x"c0",x"87",x"c4"),
  2671 => (x"4a",x"c1",x"87",x"c2"),
  2672 => (x"4f",x"26",x"48",x"72"),
  2673 => (x"4a",x"d4",x"ff",x"1e"),
  2674 => (x"c8",x"48",x"d0",x"ff"),
  2675 => (x"f0",x"c3",x"78",x"c5"),
  2676 => (x"c0",x"7a",x"71",x"7a"),
  2677 => (x"7a",x"7a",x"7a",x"7a"),
  2678 => (x"4f",x"26",x"78",x"c4"),
  2679 => (x"4a",x"d4",x"ff",x"1e"),
  2680 => (x"c8",x"48",x"d0",x"ff"),
  2681 => (x"7a",x"c0",x"78",x"c5"),
  2682 => (x"7a",x"c0",x"49",x"6a"),
  2683 => (x"7a",x"7a",x"7a",x"7a"),
  2684 => (x"48",x"71",x"78",x"c4"),
  2685 => (x"5e",x"0e",x"4f",x"26"),
  2686 => (x"0e",x"5d",x"5c",x"5b"),
  2687 => (x"a6",x"cc",x"86",x"e4"),
  2688 => (x"66",x"ec",x"c0",x"59"),
  2689 => (x"58",x"a6",x"dc",x"48"),
  2690 => (x"e4",x"c0",x"4d",x"70"),
  2691 => (x"e5",x"e4",x"c3",x"95"),
  2692 => (x"7e",x"a5",x"d4",x"85"),
  2693 => (x"d8",x"48",x"a6",x"c4"),
  2694 => (x"66",x"c4",x"78",x"a5"),
  2695 => (x"bf",x"6e",x"4c",x"bf"),
  2696 => (x"6d",x"85",x"dc",x"94"),
  2697 => (x"4b",x"66",x"c8",x"94"),
  2698 => (x"c0",x"c8",x"4a",x"c0"),
  2699 => (x"d4",x"da",x"fd",x"49"),
  2700 => (x"48",x"66",x"c8",x"87"),
  2701 => (x"78",x"9f",x"c0",x"c1"),
  2702 => (x"c2",x"49",x"66",x"c8"),
  2703 => (x"9f",x"bf",x"6e",x"81"),
  2704 => (x"49",x"66",x"c8",x"79"),
  2705 => (x"66",x"c4",x"81",x"c6"),
  2706 => (x"c8",x"79",x"9f",x"bf"),
  2707 => (x"81",x"cc",x"49",x"66"),
  2708 => (x"c8",x"79",x"9f",x"6d"),
  2709 => (x"80",x"d4",x"48",x"66"),
  2710 => (x"c2",x"58",x"a6",x"d0"),
  2711 => (x"cc",x"48",x"ec",x"ec"),
  2712 => (x"a1",x"d4",x"49",x"66"),
  2713 => (x"71",x"41",x"20",x"4a"),
  2714 => (x"87",x"f9",x"05",x"aa"),
  2715 => (x"c0",x"48",x"66",x"c8"),
  2716 => (x"a6",x"d4",x"80",x"ee"),
  2717 => (x"c1",x"ed",x"c2",x"58"),
  2718 => (x"49",x"66",x"d0",x"48"),
  2719 => (x"20",x"4a",x"a1",x"c8"),
  2720 => (x"05",x"aa",x"71",x"41"),
  2721 => (x"66",x"c8",x"87",x"f9"),
  2722 => (x"80",x"f6",x"c0",x"48"),
  2723 => (x"c2",x"58",x"a6",x"d8"),
  2724 => (x"d4",x"48",x"ca",x"ed"),
  2725 => (x"e8",x"c0",x"49",x"66"),
  2726 => (x"41",x"20",x"4a",x"a1"),
  2727 => (x"f9",x"05",x"aa",x"71"),
  2728 => (x"4a",x"66",x"d8",x"87"),
  2729 => (x"d4",x"82",x"f1",x"c0"),
  2730 => (x"81",x"cb",x"49",x"66"),
  2731 => (x"66",x"c8",x"51",x"72"),
  2732 => (x"81",x"de",x"c1",x"49"),
  2733 => (x"9f",x"d0",x"c0",x"c8"),
  2734 => (x"49",x"66",x"c8",x"79"),
  2735 => (x"c8",x"81",x"e2",x"c1"),
  2736 => (x"c8",x"79",x"9f",x"c0"),
  2737 => (x"ea",x"c1",x"49",x"66"),
  2738 => (x"79",x"9f",x"c1",x"81"),
  2739 => (x"c1",x"49",x"66",x"c8"),
  2740 => (x"bf",x"6e",x"81",x"ec"),
  2741 => (x"66",x"c8",x"79",x"9f"),
  2742 => (x"81",x"ee",x"c1",x"49"),
  2743 => (x"9f",x"bf",x"66",x"c4"),
  2744 => (x"49",x"66",x"c8",x"79"),
  2745 => (x"6d",x"81",x"f0",x"c1"),
  2746 => (x"4b",x"74",x"79",x"9f"),
  2747 => (x"9b",x"ff",x"ff",x"cf"),
  2748 => (x"66",x"c8",x"4a",x"73"),
  2749 => (x"81",x"f2",x"c1",x"49"),
  2750 => (x"74",x"79",x"9f",x"72"),
  2751 => (x"cf",x"2a",x"d0",x"4a"),
  2752 => (x"72",x"9a",x"ff",x"ff"),
  2753 => (x"49",x"66",x"c8",x"4c"),
  2754 => (x"74",x"81",x"f4",x"c1"),
  2755 => (x"c8",x"73",x"79",x"9f"),
  2756 => (x"f8",x"c1",x"49",x"66"),
  2757 => (x"79",x"9f",x"73",x"81"),
  2758 => (x"49",x"66",x"c8",x"72"),
  2759 => (x"72",x"81",x"fa",x"c1"),
  2760 => (x"8e",x"e4",x"79",x"9f"),
  2761 => (x"4c",x"26",x"4d",x"26"),
  2762 => (x"4f",x"26",x"4b",x"26"),
  2763 => (x"53",x"54",x"4d",x"69"),
  2764 => (x"6e",x"69",x"4d",x"69"),
  2765 => (x"67",x"48",x"4d",x"69"),
  2766 => (x"64",x"66",x"61",x"72"),
  2767 => (x"65",x"20",x"69",x"6c"),
  2768 => (x"30",x"31",x"2e",x"00"),
  2769 => (x"20",x"20",x"20",x"30"),
  2770 => (x"44",x"65",x"00",x"20"),
  2771 => (x"53",x"54",x"4d",x"69"),
  2772 => (x"79",x"20",x"69",x"66"),
  2773 => (x"20",x"20",x"20",x"20"),
  2774 => (x"20",x"20",x"20",x"20"),
  2775 => (x"20",x"20",x"20",x"20"),
  2776 => (x"20",x"20",x"20",x"20"),
  2777 => (x"20",x"20",x"20",x"20"),
  2778 => (x"20",x"20",x"20",x"20"),
  2779 => (x"20",x"20",x"20",x"20"),
  2780 => (x"1e",x"00",x"20",x"20"),
  2781 => (x"4b",x"71",x"1e",x"73"),
  2782 => (x"d4",x"02",x"66",x"d4"),
  2783 => (x"49",x"66",x"c8",x"87"),
  2784 => (x"4a",x"73",x"31",x"d8"),
  2785 => (x"a1",x"72",x"32",x"c8"),
  2786 => (x"81",x"66",x"cc",x"49"),
  2787 => (x"e1",x"c0",x"48",x"71"),
  2788 => (x"49",x"66",x"d0",x"87"),
  2789 => (x"c3",x"91",x"e4",x"c0"),
  2790 => (x"d8",x"81",x"e5",x"e4"),
  2791 => (x"4a",x"6a",x"4a",x"a1"),
  2792 => (x"66",x"c8",x"92",x"73"),
  2793 => (x"69",x"81",x"dc",x"82"),
  2794 => (x"cc",x"91",x"72",x"49"),
  2795 => (x"89",x"c1",x"81",x"66"),
  2796 => (x"f3",x"fd",x"48",x"71"),
  2797 => (x"4a",x"71",x"1e",x"87"),
  2798 => (x"ff",x"49",x"d4",x"ff"),
  2799 => (x"c5",x"c8",x"48",x"d0"),
  2800 => (x"79",x"d0",x"c2",x"78"),
  2801 => (x"79",x"79",x"79",x"c0"),
  2802 => (x"79",x"79",x"79",x"79"),
  2803 => (x"c0",x"79",x"72",x"79"),
  2804 => (x"79",x"66",x"c4",x"79"),
  2805 => (x"66",x"c8",x"79",x"c0"),
  2806 => (x"cc",x"79",x"c0",x"79"),
  2807 => (x"79",x"c0",x"79",x"66"),
  2808 => (x"c0",x"79",x"66",x"d0"),
  2809 => (x"79",x"66",x"d4",x"79"),
  2810 => (x"4f",x"26",x"78",x"c4"),
  2811 => (x"c6",x"4a",x"71",x"1e"),
  2812 => (x"69",x"97",x"49",x"a2"),
  2813 => (x"99",x"f0",x"c3",x"49"),
  2814 => (x"1e",x"c0",x"1e",x"71"),
  2815 => (x"c0",x"1e",x"c1",x"1e"),
  2816 => (x"f0",x"fe",x"49",x"1e"),
  2817 => (x"49",x"d0",x"c2",x"87"),
  2818 => (x"ec",x"87",x"f9",x"f6"),
  2819 => (x"1e",x"4f",x"26",x"8e"),
  2820 => (x"1e",x"1e",x"1e",x"c0"),
  2821 => (x"49",x"c1",x"1e",x"1e"),
  2822 => (x"c2",x"87",x"da",x"fe"),
  2823 => (x"e3",x"f6",x"49",x"d0"),
  2824 => (x"26",x"8e",x"ec",x"87"),
  2825 => (x"4a",x"71",x"1e",x"4f"),
  2826 => (x"c8",x"48",x"d0",x"ff"),
  2827 => (x"d4",x"ff",x"78",x"c5"),
  2828 => (x"78",x"e0",x"c2",x"48"),
  2829 => (x"78",x"78",x"78",x"c0"),
  2830 => (x"c0",x"c8",x"78",x"78"),
  2831 => (x"fd",x"49",x"72",x"1e"),
  2832 => (x"ff",x"87",x"f4",x"d3"),
  2833 => (x"78",x"c4",x"48",x"d0"),
  2834 => (x"0e",x"4f",x"26",x"26"),
  2835 => (x"5d",x"5c",x"5b",x"5e"),
  2836 => (x"71",x"86",x"f8",x"0e"),
  2837 => (x"4b",x"a2",x"c2",x"4a"),
  2838 => (x"c3",x"7b",x"97",x"c1"),
  2839 => (x"97",x"c1",x"4c",x"a2"),
  2840 => (x"c0",x"49",x"a2",x"7c"),
  2841 => (x"4d",x"a2",x"c4",x"51"),
  2842 => (x"c5",x"7d",x"97",x"c0"),
  2843 => (x"48",x"6e",x"7e",x"a2"),
  2844 => (x"a6",x"c4",x"50",x"c0"),
  2845 => (x"78",x"a2",x"c6",x"48"),
  2846 => (x"c0",x"48",x"66",x"c4"),
  2847 => (x"1e",x"66",x"d8",x"50"),
  2848 => (x"49",x"ce",x"d2",x"c3"),
  2849 => (x"c8",x"87",x"ef",x"f5"),
  2850 => (x"49",x"bf",x"97",x"66"),
  2851 => (x"97",x"66",x"c8",x"1e"),
  2852 => (x"15",x"1e",x"49",x"bf"),
  2853 => (x"49",x"14",x"1e",x"49"),
  2854 => (x"1e",x"49",x"13",x"1e"),
  2855 => (x"d4",x"fc",x"49",x"c0"),
  2856 => (x"f4",x"49",x"c8",x"87"),
  2857 => (x"d2",x"c3",x"87",x"de"),
  2858 => (x"f8",x"fd",x"49",x"ce"),
  2859 => (x"49",x"d0",x"c2",x"87"),
  2860 => (x"e0",x"87",x"d1",x"f4"),
  2861 => (x"87",x"ec",x"f9",x"8e"),
  2862 => (x"c6",x"4a",x"71",x"1e"),
  2863 => (x"69",x"97",x"49",x"a2"),
  2864 => (x"a2",x"c5",x"1e",x"49"),
  2865 => (x"49",x"69",x"97",x"49"),
  2866 => (x"49",x"a2",x"c4",x"1e"),
  2867 => (x"1e",x"49",x"69",x"97"),
  2868 => (x"97",x"49",x"a2",x"c3"),
  2869 => (x"c2",x"1e",x"49",x"69"),
  2870 => (x"69",x"97",x"49",x"a2"),
  2871 => (x"49",x"c0",x"1e",x"49"),
  2872 => (x"c2",x"87",x"d2",x"fb"),
  2873 => (x"db",x"f3",x"49",x"d0"),
  2874 => (x"26",x"8e",x"ec",x"87"),
  2875 => (x"1e",x"73",x"1e",x"4f"),
  2876 => (x"a2",x"c2",x"4a",x"71"),
  2877 => (x"d0",x"4b",x"11",x"49"),
  2878 => (x"c8",x"06",x"ab",x"b7"),
  2879 => (x"49",x"d1",x"c2",x"87"),
  2880 => (x"d5",x"87",x"c1",x"f3"),
  2881 => (x"49",x"66",x"c8",x"87"),
  2882 => (x"c3",x"91",x"e4",x"c0"),
  2883 => (x"c0",x"81",x"e5",x"e4"),
  2884 => (x"79",x"73",x"81",x"e0"),
  2885 => (x"f2",x"49",x"d0",x"c2"),
  2886 => (x"cb",x"f8",x"87",x"ea"),
  2887 => (x"1e",x"73",x"1e",x"87"),
  2888 => (x"a3",x"c6",x"4b",x"71"),
  2889 => (x"49",x"69",x"97",x"49"),
  2890 => (x"49",x"a3",x"c5",x"1e"),
  2891 => (x"1e",x"49",x"69",x"97"),
  2892 => (x"97",x"49",x"a3",x"c4"),
  2893 => (x"c3",x"1e",x"49",x"69"),
  2894 => (x"69",x"97",x"49",x"a3"),
  2895 => (x"a3",x"c2",x"1e",x"49"),
  2896 => (x"49",x"69",x"97",x"49"),
  2897 => (x"4a",x"a3",x"c1",x"1e"),
  2898 => (x"e8",x"f9",x"49",x"12"),
  2899 => (x"49",x"d0",x"c2",x"87"),
  2900 => (x"ec",x"87",x"f1",x"f1"),
  2901 => (x"87",x"d0",x"f7",x"8e"),
  2902 => (x"5c",x"5b",x"5e",x"0e"),
  2903 => (x"71",x"1e",x"0e",x"5d"),
  2904 => (x"c2",x"49",x"6e",x"7e"),
  2905 => (x"79",x"97",x"c1",x"81"),
  2906 => (x"83",x"c3",x"4b",x"6e"),
  2907 => (x"6e",x"7b",x"97",x"c1"),
  2908 => (x"c0",x"82",x"c1",x"4a"),
  2909 => (x"4c",x"6e",x"7a",x"97"),
  2910 => (x"97",x"c0",x"84",x"c4"),
  2911 => (x"c5",x"4d",x"6e",x"7c"),
  2912 => (x"6e",x"55",x"c0",x"85"),
  2913 => (x"97",x"85",x"c6",x"4d"),
  2914 => (x"c0",x"1e",x"4d",x"6d"),
  2915 => (x"4c",x"6c",x"97",x"1e"),
  2916 => (x"4b",x"6b",x"97",x"1e"),
  2917 => (x"49",x"69",x"97",x"1e"),
  2918 => (x"f8",x"49",x"12",x"1e"),
  2919 => (x"d0",x"c2",x"87",x"d7"),
  2920 => (x"87",x"e0",x"f0",x"49"),
  2921 => (x"fb",x"f5",x"8e",x"e8"),
  2922 => (x"5b",x"5e",x"0e",x"87"),
  2923 => (x"ff",x"0e",x"5d",x"5c"),
  2924 => (x"4b",x"71",x"86",x"dc"),
  2925 => (x"11",x"49",x"a3",x"c3"),
  2926 => (x"58",x"a6",x"d4",x"48"),
  2927 => (x"c5",x"4a",x"a3",x"c4"),
  2928 => (x"69",x"97",x"49",x"a3"),
  2929 => (x"97",x"31",x"c8",x"49"),
  2930 => (x"71",x"48",x"4a",x"6a"),
  2931 => (x"58",x"a6",x"d8",x"b0"),
  2932 => (x"6e",x"7e",x"a3",x"c6"),
  2933 => (x"4d",x"49",x"bf",x"97"),
  2934 => (x"48",x"71",x"9d",x"cf"),
  2935 => (x"dc",x"98",x"c0",x"c1"),
  2936 => (x"ec",x"48",x"58",x"a6"),
  2937 => (x"78",x"a3",x"c2",x"80"),
  2938 => (x"bf",x"97",x"66",x"c4"),
  2939 => (x"c3",x"05",x"9c",x"4c"),
  2940 => (x"4c",x"c0",x"c4",x"87"),
  2941 => (x"c0",x"1e",x"66",x"d8"),
  2942 => (x"d8",x"1e",x"66",x"f8"),
  2943 => (x"1e",x"75",x"1e",x"66"),
  2944 => (x"49",x"66",x"e4",x"c0"),
  2945 => (x"d0",x"87",x"ec",x"f5"),
  2946 => (x"c0",x"49",x"70",x"86"),
  2947 => (x"74",x"59",x"a6",x"e0"),
  2948 => (x"fb",x"c5",x"02",x"9c"),
  2949 => (x"66",x"f8",x"c0",x"87"),
  2950 => (x"d0",x"87",x"c5",x"02"),
  2951 => (x"87",x"c5",x"5c",x"a6"),
  2952 => (x"c1",x"48",x"a6",x"cc"),
  2953 => (x"4b",x"66",x"cc",x"78"),
  2954 => (x"02",x"66",x"f8",x"c0"),
  2955 => (x"f4",x"c0",x"87",x"de"),
  2956 => (x"e4",x"c0",x"49",x"66"),
  2957 => (x"e5",x"e4",x"c3",x"91"),
  2958 => (x"81",x"e0",x"c0",x"81"),
  2959 => (x"69",x"48",x"a6",x"c8"),
  2960 => (x"48",x"66",x"cc",x"78"),
  2961 => (x"a8",x"b7",x"66",x"c8"),
  2962 => (x"4b",x"87",x"c1",x"06"),
  2963 => (x"05",x"66",x"fc",x"c0"),
  2964 => (x"49",x"c8",x"87",x"d9"),
  2965 => (x"ee",x"87",x"ed",x"ed"),
  2966 => (x"49",x"70",x"87",x"c2"),
  2967 => (x"ca",x"05",x"99",x"c4"),
  2968 => (x"87",x"f8",x"ed",x"87"),
  2969 => (x"99",x"c4",x"49",x"70"),
  2970 => (x"73",x"87",x"f6",x"02"),
  2971 => (x"d0",x"88",x"c1",x"48"),
  2972 => (x"4a",x"70",x"58",x"a6"),
  2973 => (x"c1",x"02",x"9b",x"73"),
  2974 => (x"ac",x"c1",x"87",x"d3"),
  2975 => (x"87",x"c1",x"c1",x"02"),
  2976 => (x"49",x"66",x"f4",x"c0"),
  2977 => (x"c3",x"91",x"e4",x"c0"),
  2978 => (x"71",x"48",x"e5",x"e4"),
  2979 => (x"58",x"a6",x"cc",x"80"),
  2980 => (x"dc",x"49",x"66",x"c8"),
  2981 => (x"48",x"66",x"d0",x"81"),
  2982 => (x"dc",x"05",x"a8",x"69"),
  2983 => (x"48",x"a6",x"d0",x"87"),
  2984 => (x"c8",x"85",x"78",x"c1"),
  2985 => (x"81",x"d8",x"49",x"66"),
  2986 => (x"d4",x"05",x"ad",x"69"),
  2987 => (x"d4",x"4d",x"c0",x"87"),
  2988 => (x"80",x"c1",x"48",x"66"),
  2989 => (x"c8",x"58",x"a6",x"d8"),
  2990 => (x"48",x"66",x"d0",x"87"),
  2991 => (x"a6",x"d4",x"80",x"c1"),
  2992 => (x"72",x"8c",x"c1",x"58"),
  2993 => (x"71",x"8a",x"c1",x"49"),
  2994 => (x"ed",x"fe",x"05",x"99"),
  2995 => (x"02",x"66",x"d8",x"87"),
  2996 => (x"49",x"73",x"87",x"da"),
  2997 => (x"71",x"81",x"66",x"dc"),
  2998 => (x"9a",x"ff",x"c3",x"4a"),
  2999 => (x"71",x"5a",x"a6",x"d4"),
  3000 => (x"2a",x"b7",x"c8",x"4a"),
  3001 => (x"d8",x"5a",x"a6",x"d8"),
  3002 => (x"4d",x"71",x"29",x"b7"),
  3003 => (x"49",x"bf",x"97",x"6e"),
  3004 => (x"75",x"99",x"f0",x"c3"),
  3005 => (x"d8",x"1e",x"71",x"b1"),
  3006 => (x"b7",x"c8",x"49",x"66"),
  3007 => (x"dc",x"1e",x"71",x"29"),
  3008 => (x"66",x"dc",x"1e",x"66"),
  3009 => (x"97",x"66",x"d4",x"1e"),
  3010 => (x"c0",x"1e",x"49",x"bf"),
  3011 => (x"87",x"e5",x"f2",x"49"),
  3012 => (x"fc",x"c0",x"86",x"d4"),
  3013 => (x"f1",x"c1",x"05",x"66"),
  3014 => (x"ea",x"49",x"d0",x"87"),
  3015 => (x"f4",x"c0",x"87",x"e6"),
  3016 => (x"e4",x"c0",x"49",x"66"),
  3017 => (x"e5",x"e4",x"c3",x"91"),
  3018 => (x"cc",x"80",x"71",x"48"),
  3019 => (x"66",x"c8",x"58",x"a6"),
  3020 => (x"69",x"81",x"c8",x"49"),
  3021 => (x"87",x"cd",x"c1",x"02"),
  3022 => (x"c9",x"49",x"66",x"dc"),
  3023 => (x"cc",x"1e",x"71",x"31"),
  3024 => (x"ec",x"fd",x"49",x"66"),
  3025 => (x"86",x"c4",x"87",x"ce"),
  3026 => (x"48",x"a6",x"e0",x"c0"),
  3027 => (x"73",x"78",x"66",x"cc"),
  3028 => (x"f5",x"c0",x"02",x"9b"),
  3029 => (x"cc",x"1e",x"c0",x"87"),
  3030 => (x"e9",x"fd",x"49",x"66"),
  3031 => (x"1e",x"c1",x"87",x"d8"),
  3032 => (x"fd",x"49",x"66",x"d0"),
  3033 => (x"c8",x"87",x"f5",x"e7"),
  3034 => (x"48",x"66",x"dc",x"86"),
  3035 => (x"e0",x"c0",x"80",x"c1"),
  3036 => (x"e0",x"c0",x"58",x"a6"),
  3037 => (x"c1",x"48",x"49",x"66"),
  3038 => (x"a6",x"e4",x"c0",x"88"),
  3039 => (x"05",x"99",x"71",x"58"),
  3040 => (x"c5",x"87",x"d2",x"ff"),
  3041 => (x"e8",x"49",x"c9",x"87"),
  3042 => (x"9c",x"74",x"87",x"fa"),
  3043 => (x"87",x"c5",x"fa",x"05"),
  3044 => (x"02",x"66",x"fc",x"c0"),
  3045 => (x"d0",x"c2",x"87",x"c8"),
  3046 => (x"87",x"e8",x"e8",x"49"),
  3047 => (x"c0",x"c2",x"87",x"c6"),
  3048 => (x"87",x"e0",x"e8",x"49"),
  3049 => (x"ed",x"8e",x"dc",x"ff"),
  3050 => (x"5e",x"0e",x"87",x"fa"),
  3051 => (x"0e",x"5d",x"5c",x"5b"),
  3052 => (x"4c",x"71",x"86",x"e0"),
  3053 => (x"11",x"49",x"a4",x"c3"),
  3054 => (x"58",x"a6",x"d4",x"48"),
  3055 => (x"c5",x"4a",x"a4",x"c4"),
  3056 => (x"69",x"97",x"49",x"a4"),
  3057 => (x"97",x"31",x"c8",x"49"),
  3058 => (x"71",x"48",x"4a",x"6a"),
  3059 => (x"58",x"a6",x"d8",x"b0"),
  3060 => (x"6e",x"7e",x"a4",x"c6"),
  3061 => (x"4d",x"49",x"bf",x"97"),
  3062 => (x"48",x"71",x"9d",x"cf"),
  3063 => (x"dc",x"98",x"c0",x"c1"),
  3064 => (x"ec",x"48",x"58",x"a6"),
  3065 => (x"78",x"a4",x"c2",x"80"),
  3066 => (x"bf",x"97",x"66",x"c4"),
  3067 => (x"1e",x"66",x"d8",x"4b"),
  3068 => (x"1e",x"66",x"f4",x"c0"),
  3069 => (x"75",x"1e",x"66",x"d8"),
  3070 => (x"66",x"e4",x"c0",x"1e"),
  3071 => (x"87",x"f3",x"ed",x"49"),
  3072 => (x"49",x"70",x"86",x"d0"),
  3073 => (x"59",x"a6",x"e0",x"c0"),
  3074 => (x"c3",x"05",x"9b",x"73"),
  3075 => (x"4b",x"c0",x"c4",x"87"),
  3076 => (x"ef",x"e6",x"49",x"c4"),
  3077 => (x"49",x"66",x"dc",x"87"),
  3078 => (x"1e",x"71",x"31",x"c9"),
  3079 => (x"49",x"66",x"f4",x"c0"),
  3080 => (x"c3",x"91",x"e4",x"c0"),
  3081 => (x"71",x"48",x"e5",x"e4"),
  3082 => (x"58",x"a6",x"d4",x"80"),
  3083 => (x"fd",x"49",x"66",x"d0"),
  3084 => (x"c4",x"87",x"e1",x"e8"),
  3085 => (x"02",x"9b",x"73",x"86"),
  3086 => (x"c0",x"87",x"dd",x"c4"),
  3087 => (x"c4",x"02",x"66",x"f4"),
  3088 => (x"c2",x"4a",x"73",x"87"),
  3089 => (x"72",x"4a",x"c1",x"87"),
  3090 => (x"66",x"f4",x"c0",x"4c"),
  3091 => (x"cc",x"87",x"d3",x"02"),
  3092 => (x"e0",x"c0",x"49",x"66"),
  3093 => (x"48",x"a6",x"c8",x"81"),
  3094 => (x"66",x"c8",x"78",x"69"),
  3095 => (x"c1",x"06",x"aa",x"b7"),
  3096 => (x"9c",x"74",x"4c",x"87"),
  3097 => (x"87",x"d3",x"c2",x"02"),
  3098 => (x"70",x"87",x"f1",x"e5"),
  3099 => (x"05",x"99",x"c8",x"49"),
  3100 => (x"e7",x"e5",x"87",x"ca"),
  3101 => (x"c8",x"49",x"70",x"87"),
  3102 => (x"87",x"f6",x"02",x"99"),
  3103 => (x"c8",x"48",x"d0",x"ff"),
  3104 => (x"d4",x"ff",x"78",x"c5"),
  3105 => (x"78",x"f0",x"c2",x"48"),
  3106 => (x"78",x"78",x"78",x"c0"),
  3107 => (x"c0",x"c8",x"78",x"78"),
  3108 => (x"ce",x"d2",x"c3",x"1e"),
  3109 => (x"c5",x"c3",x"fd",x"49"),
  3110 => (x"48",x"d0",x"ff",x"87"),
  3111 => (x"d2",x"c3",x"78",x"c4"),
  3112 => (x"66",x"d4",x"1e",x"ce"),
  3113 => (x"dc",x"e5",x"fd",x"49"),
  3114 => (x"d8",x"1e",x"c1",x"87"),
  3115 => (x"e2",x"fd",x"49",x"66"),
  3116 => (x"86",x"cc",x"87",x"ea"),
  3117 => (x"c1",x"48",x"66",x"dc"),
  3118 => (x"a6",x"e0",x"c0",x"80"),
  3119 => (x"02",x"ab",x"c1",x"58"),
  3120 => (x"cc",x"87",x"f1",x"c0"),
  3121 => (x"81",x"dc",x"49",x"66"),
  3122 => (x"69",x"48",x"66",x"d0"),
  3123 => (x"87",x"dc",x"05",x"a8"),
  3124 => (x"c1",x"48",x"a6",x"d0"),
  3125 => (x"66",x"cc",x"85",x"78"),
  3126 => (x"69",x"81",x"d8",x"49"),
  3127 => (x"87",x"d4",x"05",x"ad"),
  3128 => (x"66",x"d4",x"4d",x"c0"),
  3129 => (x"d8",x"80",x"c1",x"48"),
  3130 => (x"87",x"c8",x"58",x"a6"),
  3131 => (x"c1",x"48",x"66",x"d0"),
  3132 => (x"58",x"a6",x"d4",x"80"),
  3133 => (x"05",x"8c",x"8b",x"c1"),
  3134 => (x"d8",x"87",x"ed",x"fd"),
  3135 => (x"87",x"da",x"02",x"66"),
  3136 => (x"c3",x"49",x"66",x"dc"),
  3137 => (x"a6",x"d4",x"99",x"ff"),
  3138 => (x"49",x"66",x"dc",x"59"),
  3139 => (x"d8",x"29",x"b7",x"c8"),
  3140 => (x"66",x"dc",x"59",x"a6"),
  3141 => (x"29",x"b7",x"d8",x"49"),
  3142 => (x"97",x"6e",x"4d",x"71"),
  3143 => (x"f0",x"c3",x"49",x"bf"),
  3144 => (x"71",x"b1",x"75",x"99"),
  3145 => (x"49",x"66",x"d8",x"1e"),
  3146 => (x"71",x"29",x"b7",x"c8"),
  3147 => (x"1e",x"66",x"dc",x"1e"),
  3148 => (x"d4",x"1e",x"66",x"dc"),
  3149 => (x"49",x"bf",x"97",x"66"),
  3150 => (x"e9",x"49",x"c0",x"1e"),
  3151 => (x"86",x"d4",x"87",x"f7"),
  3152 => (x"c7",x"02",x"9b",x"73"),
  3153 => (x"e1",x"49",x"d0",x"87"),
  3154 => (x"87",x"c6",x"87",x"fa"),
  3155 => (x"e1",x"49",x"d0",x"c2"),
  3156 => (x"9b",x"73",x"87",x"f2"),
  3157 => (x"87",x"e3",x"fb",x"05"),
  3158 => (x"c7",x"e7",x"8e",x"e0"),
  3159 => (x"5b",x"5e",x"0e",x"87"),
  3160 => (x"e4",x"0e",x"5d",x"5c"),
  3161 => (x"cc",x"4a",x"71",x"86"),
  3162 => (x"ff",x"c0",x"48",x"a6"),
  3163 => (x"c1",x"80",x"c4",x"78"),
  3164 => (x"80",x"c4",x"78",x"ff"),
  3165 => (x"c4",x"78",x"ff",x"c3"),
  3166 => (x"c8",x"78",x"c0",x"80"),
  3167 => (x"49",x"69",x"49",x"a2"),
  3168 => (x"4d",x"71",x"29",x"c9"),
  3169 => (x"eb",x"c2",x"02",x"9d"),
  3170 => (x"cc",x"4c",x"c0",x"87"),
  3171 => (x"02",x"6b",x"4b",x"a6"),
  3172 => (x"74",x"87",x"ca",x"c2"),
  3173 => (x"73",x"91",x"c4",x"49"),
  3174 => (x"7e",x"69",x"49",x"a1"),
  3175 => (x"c4",x"48",x"a6",x"c8"),
  3176 => (x"49",x"66",x"c8",x"78"),
  3177 => (x"1e",x"71",x"91",x"6e"),
  3178 => (x"09",x"75",x"1e",x"72"),
  3179 => (x"d5",x"fd",x"fc",x"4a"),
  3180 => (x"26",x"4a",x"26",x"87"),
  3181 => (x"58",x"a6",x"c8",x"49"),
  3182 => (x"c0",x"c0",x"c0",x"c4"),
  3183 => (x"cb",x"01",x"ad",x"b7"),
  3184 => (x"b7",x"ff",x"cf",x"87"),
  3185 => (x"fd",x"c0",x"06",x"a8"),
  3186 => (x"87",x"eb",x"c0",x"87"),
  3187 => (x"c3",x"48",x"66",x"c4"),
  3188 => (x"a8",x"b7",x"ff",x"ff"),
  3189 => (x"87",x"ee",x"c0",x"04"),
  3190 => (x"c7",x"48",x"66",x"c4"),
  3191 => (x"a8",x"b7",x"ff",x"ff"),
  3192 => (x"c8",x"87",x"c9",x"03"),
  3193 => (x"b7",x"c5",x"48",x"66"),
  3194 => (x"87",x"da",x"03",x"a8"),
  3195 => (x"cf",x"48",x"66",x"c4"),
  3196 => (x"a8",x"b7",x"ff",x"ff"),
  3197 => (x"c8",x"87",x"cf",x"06"),
  3198 => (x"80",x"c1",x"48",x"66"),
  3199 => (x"d0",x"58",x"a6",x"cc"),
  3200 => (x"fe",x"06",x"a8",x"b7"),
  3201 => (x"66",x"c8",x"87",x"db"),
  3202 => (x"a8",x"b7",x"d0",x"48"),
  3203 => (x"c1",x"87",x"ce",x"06"),
  3204 => (x"c4",x"49",x"74",x"84"),
  3205 => (x"49",x"a1",x"73",x"91"),
  3206 => (x"f6",x"fd",x"05",x"69"),
  3207 => (x"49",x"a2",x"d4",x"87"),
  3208 => (x"d8",x"79",x"66",x"c4"),
  3209 => (x"66",x"c8",x"49",x"a2"),
  3210 => (x"49",x"a2",x"dc",x"79"),
  3211 => (x"e0",x"c0",x"79",x"6e"),
  3212 => (x"79",x"c1",x"49",x"a2"),
  3213 => (x"eb",x"e3",x"8e",x"e4"),
  3214 => (x"49",x"c0",x"1e",x"87"),
  3215 => (x"bf",x"ed",x"e4",x"c3"),
  3216 => (x"c1",x"87",x"c2",x"02"),
  3217 => (x"d1",x"e5",x"c3",x"49"),
  3218 => (x"87",x"c2",x"02",x"bf"),
  3219 => (x"d0",x"ff",x"b1",x"c2"),
  3220 => (x"78",x"c5",x"c8",x"48"),
  3221 => (x"c3",x"48",x"d4",x"ff"),
  3222 => (x"78",x"71",x"78",x"fa"),
  3223 => (x"c4",x"48",x"d0",x"ff"),
  3224 => (x"1e",x"4f",x"26",x"78"),
  3225 => (x"4a",x"71",x"1e",x"73"),
  3226 => (x"49",x"66",x"cc",x"1e"),
  3227 => (x"c3",x"91",x"e4",x"c0"),
  3228 => (x"71",x"4b",x"e5",x"e4"),
  3229 => (x"fd",x"49",x"73",x"83"),
  3230 => (x"c4",x"87",x"e6",x"d9"),
  3231 => (x"02",x"98",x"70",x"86"),
  3232 => (x"49",x"73",x"87",x"c5"),
  3233 => (x"fe",x"87",x"d6",x"fb"),
  3234 => (x"db",x"e2",x"87",x"ef"),
  3235 => (x"5b",x"5e",x"0e",x"87"),
  3236 => (x"f4",x"0e",x"5d",x"5c"),
  3237 => (x"c3",x"dd",x"ff",x"86"),
  3238 => (x"c4",x"49",x"70",x"87"),
  3239 => (x"ec",x"c5",x"02",x"99"),
  3240 => (x"48",x"d0",x"ff",x"87"),
  3241 => (x"ff",x"78",x"c5",x"c8"),
  3242 => (x"c0",x"c2",x"48",x"d4"),
  3243 => (x"78",x"78",x"c0",x"78"),
  3244 => (x"4d",x"78",x"78",x"78"),
  3245 => (x"c0",x"48",x"d4",x"ff"),
  3246 => (x"a5",x"4a",x"76",x"78"),
  3247 => (x"bf",x"d4",x"ff",x"49"),
  3248 => (x"d4",x"ff",x"79",x"97"),
  3249 => (x"68",x"78",x"c0",x"48"),
  3250 => (x"c8",x"85",x"c1",x"51"),
  3251 => (x"e3",x"04",x"ad",x"b7"),
  3252 => (x"48",x"d0",x"ff",x"87"),
  3253 => (x"97",x"c6",x"78",x"c4"),
  3254 => (x"a6",x"cc",x"48",x"66"),
  3255 => (x"d0",x"4b",x"70",x"58"),
  3256 => (x"2b",x"b7",x"c4",x"9b"),
  3257 => (x"e4",x"c0",x"49",x"73"),
  3258 => (x"e5",x"e4",x"c3",x"91"),
  3259 => (x"69",x"81",x"c8",x"81"),
  3260 => (x"c2",x"87",x"ca",x"05"),
  3261 => (x"db",x"ff",x"49",x"d1"),
  3262 => (x"d0",x"c4",x"87",x"ca"),
  3263 => (x"66",x"97",x"c7",x"87"),
  3264 => (x"f0",x"c3",x"49",x"4c"),
  3265 => (x"05",x"a9",x"d0",x"99"),
  3266 => (x"1e",x"73",x"87",x"cc"),
  3267 => (x"db",x"e3",x"49",x"72"),
  3268 => (x"c3",x"86",x"c4",x"87"),
  3269 => (x"d0",x"c2",x"87",x"f7"),
  3270 => (x"87",x"c8",x"05",x"ac"),
  3271 => (x"ee",x"e3",x"49",x"72"),
  3272 => (x"87",x"e9",x"c3",x"87"),
  3273 => (x"05",x"ac",x"ec",x"c3"),
  3274 => (x"1e",x"c0",x"87",x"ce"),
  3275 => (x"49",x"72",x"1e",x"73"),
  3276 => (x"c8",x"87",x"d8",x"e4"),
  3277 => (x"87",x"d5",x"c3",x"86"),
  3278 => (x"05",x"ac",x"d1",x"c2"),
  3279 => (x"1e",x"73",x"87",x"cc"),
  3280 => (x"f3",x"e5",x"49",x"72"),
  3281 => (x"c3",x"86",x"c4",x"87"),
  3282 => (x"c6",x"c3",x"87",x"c3"),
  3283 => (x"87",x"cc",x"05",x"ac"),
  3284 => (x"49",x"72",x"1e",x"73"),
  3285 => (x"c4",x"87",x"d6",x"e6"),
  3286 => (x"87",x"f1",x"c2",x"86"),
  3287 => (x"05",x"ac",x"e0",x"c0"),
  3288 => (x"1e",x"c0",x"87",x"cf"),
  3289 => (x"72",x"1e",x"73",x"1e"),
  3290 => (x"87",x"fd",x"e8",x"49"),
  3291 => (x"dc",x"c2",x"86",x"cc"),
  3292 => (x"ac",x"c4",x"c3",x"87"),
  3293 => (x"c0",x"87",x"d0",x"05"),
  3294 => (x"73",x"1e",x"c1",x"1e"),
  3295 => (x"e8",x"49",x"72",x"1e"),
  3296 => (x"86",x"cc",x"87",x"e7"),
  3297 => (x"c0",x"87",x"c6",x"c2"),
  3298 => (x"ce",x"05",x"ac",x"f0"),
  3299 => (x"73",x"1e",x"c0",x"87"),
  3300 => (x"f0",x"49",x"72",x"1e"),
  3301 => (x"86",x"c8",x"87",x"d4"),
  3302 => (x"c3",x"87",x"f2",x"c1"),
  3303 => (x"ce",x"05",x"ac",x"c5"),
  3304 => (x"73",x"1e",x"c1",x"87"),
  3305 => (x"f0",x"49",x"72",x"1e"),
  3306 => (x"86",x"c8",x"87",x"c0"),
  3307 => (x"c8",x"87",x"de",x"c1"),
  3308 => (x"87",x"cc",x"05",x"ac"),
  3309 => (x"49",x"72",x"1e",x"73"),
  3310 => (x"c4",x"87",x"dd",x"e6"),
  3311 => (x"87",x"cd",x"c1",x"86"),
  3312 => (x"05",x"ac",x"c0",x"c1"),
  3313 => (x"1e",x"c1",x"87",x"d0"),
  3314 => (x"1e",x"73",x"1e",x"c0"),
  3315 => (x"d8",x"e7",x"49",x"72"),
  3316 => (x"c0",x"86",x"cc",x"87"),
  3317 => (x"9c",x"74",x"87",x"f7"),
  3318 => (x"73",x"87",x"cc",x"05"),
  3319 => (x"e4",x"49",x"72",x"1e"),
  3320 => (x"86",x"c4",x"87",x"fb"),
  3321 => (x"c8",x"87",x"e6",x"c0"),
  3322 => (x"97",x"c9",x"1e",x"66"),
  3323 => (x"cc",x"1e",x"49",x"66"),
  3324 => (x"1e",x"49",x"66",x"97"),
  3325 => (x"49",x"66",x"97",x"cf"),
  3326 => (x"66",x"97",x"d2",x"1e"),
  3327 => (x"49",x"c4",x"1e",x"49"),
  3328 => (x"87",x"f1",x"de",x"ff"),
  3329 => (x"d1",x"c2",x"86",x"d4"),
  3330 => (x"f7",x"d6",x"ff",x"49"),
  3331 => (x"ff",x"8e",x"f4",x"87"),
  3332 => (x"1e",x"87",x"d1",x"dc"),
  3333 => (x"bf",x"e1",x"d1",x"c3"),
  3334 => (x"c3",x"b9",x"c1",x"49"),
  3335 => (x"ff",x"59",x"e5",x"d1"),
  3336 => (x"ff",x"c3",x"48",x"d4"),
  3337 => (x"48",x"d0",x"ff",x"78"),
  3338 => (x"ff",x"78",x"e1",x"c8"),
  3339 => (x"78",x"c1",x"48",x"d4"),
  3340 => (x"78",x"71",x"31",x"c4"),
  3341 => (x"c0",x"48",x"d0",x"ff"),
  3342 => (x"4f",x"26",x"78",x"e0"),
  3343 => (x"d5",x"d1",x"c3",x"1e"),
  3344 => (x"c4",x"df",x"c3",x"1e"),
  3345 => (x"d8",x"d2",x"fd",x"49"),
  3346 => (x"70",x"86",x"c4",x"87"),
  3347 => (x"87",x"c3",x"02",x"98"),
  3348 => (x"26",x"87",x"c0",x"ff"),
  3349 => (x"4b",x"35",x"31",x"4f"),
  3350 => (x"20",x"20",x"5a",x"48"),
  3351 => (x"47",x"46",x"43",x"20"),
  3352 => (x"00",x"00",x"00",x"00"),
  3353 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

