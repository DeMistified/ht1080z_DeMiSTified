library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"486e87c4",
     1 => x"66c850c0",
     2 => x"c387c705",
     3 => x"c448e4e3",
     4 => x"85c178a5",
     5 => x"04adb7c4",
     6 => x"c487c0ff",
     7 => x"e3c387dc",
     8 => x"c848bff0",
     9 => x"d101a8b7",
    10 => x"02acca87",
    11 => x"accd87cc",
    12 => x"c087c702",
    13 => x"c003acb7",
    14 => x"e3c387f3",
    15 => x"c84bbff0",
    16 => x"d203abb7",
    17 => x"f4e3c387",
    18 => x"c0817349",
    19 => x"83c151e0",
    20 => x"04abb7c8",
    21 => x"c387eeff",
    22 => x"c148fce3",
    23 => x"cfc150d2",
    24 => x"50cdc150",
    25 => x"80e450c0",
    26 => x"cdc378c3",
    27 => x"f0e3c387",
    28 => x"c14849bf",
    29 => x"f4e3c380",
    30 => x"a0c44858",
    31 => x"c2517481",
    32 => x"f0c087f8",
    33 => x"da04acb7",
    34 => x"b7f9c087",
    35 => x"87d301ac",
    36 => x"bfe8e3c3",
    37 => x"7491ca49",
    38 => x"8af0c04a",
    39 => x"48e8e3c3",
    40 => x"ca78a172",
    41 => x"c6c002ac",
    42 => x"05accd87",
    43 => x"c387cbc2",
    44 => x"c348e4e3",
    45 => x"87c2c278",
    46 => x"acb7f0c0",
    47 => x"c087db04",
    48 => x"01acb7f9",
    49 => x"c387d3c0",
    50 => x"49bfece3",
    51 => x"4a7491d0",
    52 => x"c38af0c0",
    53 => x"7248ece3",
    54 => x"c1c178a1",
    55 => x"c004acb7",
    56 => x"c6c187db",
    57 => x"c001acb7",
    58 => x"e3c387d3",
    59 => x"d049bfec",
    60 => x"c04a7491",
    61 => x"e3c38af7",
    62 => x"a17248ec",
    63 => x"02acca78",
    64 => x"cd87c6c0",
    65 => x"f1c005ac",
    66 => x"e4e3c387",
    67 => x"c078c348",
    68 => x"e2c087e8",
    69 => x"c9c005ac",
    70 => x"48a6c487",
    71 => x"c078fbc0",
    72 => x"acca87d8",
    73 => x"87c6c002",
    74 => x"c005accd",
    75 => x"e3c387c9",
    76 => x"78c348e4",
    77 => x"c887c3c0",
    78 => x"b7c05ca6",
    79 => x"c4c003ac",
    80 => x"cac04887",
    81 => x"0266c487",
    82 => x"4887c6f9",
    83 => x"f499ffc3",
    84 => x"87cff88e",
    85 => x"464e4f43",
    86 => x"4f4d003d",
    87 => x"414e0044",
    88 => x"4400454d",
    89 => x"55414645",
    90 => x"303d544c",
    91 => x"00215400",
    92 => x"00215a00",
    93 => x"00215e00",
    94 => x"00216300",
    95 => x"d0ff1e00",
    96 => x"78c9c848",
    97 => x"d4ff4871",
    98 => x"4f267808",
    99 => x"494a711e",
   100 => x"d0ff87eb",
   101 => x"2678c848",
   102 => x"1e731e4f",
   103 => x"e4c34b71",
   104 => x"c302bfcc",
   105 => x"87ebc287",
   106 => x"c848d0ff",
   107 => x"497378c9",
   108 => x"ffb1e0c0",
   109 => x"787148d4",
   110 => x"48c0e4c3",
   111 => x"66c878c0",
   112 => x"c387c502",
   113 => x"87c249ff",
   114 => x"e4c349c0",
   115 => x"66cc59c8",
   116 => x"c587c602",
   117 => x"c44ad5d5",
   118 => x"ffffcf87",
   119 => x"cce4c34a",
   120 => x"cce4c35a",
   121 => x"c478c148",
   122 => x"264d2687",
   123 => x"264b264c",
   124 => x"5b5e0e4f",
   125 => x"710e5d5c",
   126 => x"c8e4c34a",
   127 => x"9a724cbf",
   128 => x"4987cb02",
   129 => x"c6c291c8",
   130 => x"83714bcf",
   131 => x"cac287c4",
   132 => x"4dc04bcf",
   133 => x"99744913",
   134 => x"bfc4e4c3",
   135 => x"48d4ffb9",
   136 => x"b7c17871",
   137 => x"b7c8852c",
   138 => x"87e804ad",
   139 => x"bfc0e4c3",
   140 => x"c380c848",
   141 => x"fe58c4e4",
   142 => x"731e87ef",
   143 => x"134b711e",
   144 => x"cb029a4a",
   145 => x"fe497287",
   146 => x"4a1387e7",
   147 => x"87f5059a",
   148 => x"1e87dafe",
   149 => x"bfc0e4c3",
   150 => x"c0e4c349",
   151 => x"78a1c148",
   152 => x"a9b7c0c4",
   153 => x"ff87db03",
   154 => x"e4c348d4",
   155 => x"c378bfc4",
   156 => x"49bfc0e4",
   157 => x"48c0e4c3",
   158 => x"c478a1c1",
   159 => x"04a9b7c0",
   160 => x"d0ff87e5",
   161 => x"c378c848",
   162 => x"c048cce4",
   163 => x"004f2678",
   164 => x"00000000",
   165 => x"00000000",
   166 => x"5f5f0000",
   167 => x"00000000",
   168 => x"03000303",
   169 => x"14000003",
   170 => x"7f147f7f",
   171 => x"0000147f",
   172 => x"6b6b2e24",
   173 => x"4c00123a",
   174 => x"6c18366a",
   175 => x"30003256",
   176 => x"77594f7e",
   177 => x"0040683a",
   178 => x"03070400",
   179 => x"00000000",
   180 => x"633e1c00",
   181 => x"00000041",
   182 => x"3e634100",
   183 => x"0800001c",
   184 => x"1c1c3e2a",
   185 => x"00082a3e",
   186 => x"3e3e0808",
   187 => x"00000808",
   188 => x"60e08000",
   189 => x"00000000",
   190 => x"08080808",
   191 => x"00000808",
   192 => x"60600000",
   193 => x"40000000",
   194 => x"0c183060",
   195 => x"00010306",
   196 => x"4d597f3e",
   197 => x"00003e7f",
   198 => x"7f7f0604",
   199 => x"00000000",
   200 => x"59716342",
   201 => x"0000464f",
   202 => x"49496322",
   203 => x"1800367f",
   204 => x"7f13161c",
   205 => x"0000107f",
   206 => x"45456727",
   207 => x"0000397d",
   208 => x"494b7e3c",
   209 => x"00003079",
   210 => x"79710101",
   211 => x"0000070f",
   212 => x"49497f36",
   213 => x"0000367f",
   214 => x"69494f06",
   215 => x"00001e3f",
   216 => x"66660000",
   217 => x"00000000",
   218 => x"66e68000",
   219 => x"00000000",
   220 => x"14140808",
   221 => x"00002222",
   222 => x"14141414",
   223 => x"00001414",
   224 => x"14142222",
   225 => x"00000808",
   226 => x"59510302",
   227 => x"3e00060f",
   228 => x"555d417f",
   229 => x"00001e1f",
   230 => x"09097f7e",
   231 => x"00007e7f",
   232 => x"49497f7f",
   233 => x"0000367f",
   234 => x"41633e1c",
   235 => x"00004141",
   236 => x"63417f7f",
   237 => x"00001c3e",
   238 => x"49497f7f",
   239 => x"00004141",
   240 => x"09097f7f",
   241 => x"00000101",
   242 => x"49417f3e",
   243 => x"00007a7b",
   244 => x"08087f7f",
   245 => x"00007f7f",
   246 => x"7f7f4100",
   247 => x"00000041",
   248 => x"40406020",
   249 => x"7f003f7f",
   250 => x"361c087f",
   251 => x"00004163",
   252 => x"40407f7f",
   253 => x"7f004040",
   254 => x"060c067f",
   255 => x"7f007f7f",
   256 => x"180c067f",
   257 => x"00007f7f",
   258 => x"41417f3e",
   259 => x"00003e7f",
   260 => x"09097f7f",
   261 => x"3e00060f",
   262 => x"7f61417f",
   263 => x"0000407e",
   264 => x"19097f7f",
   265 => x"0000667f",
   266 => x"594d6f26",
   267 => x"0000327b",
   268 => x"7f7f0101",
   269 => x"00000101",
   270 => x"40407f3f",
   271 => x"00003f7f",
   272 => x"70703f0f",
   273 => x"7f000f3f",
   274 => x"3018307f",
   275 => x"41007f7f",
   276 => x"1c1c3663",
   277 => x"01416336",
   278 => x"7c7c0603",
   279 => x"61010306",
   280 => x"474d5971",
   281 => x"00004143",
   282 => x"417f7f00",
   283 => x"01000041",
   284 => x"180c0603",
   285 => x"00406030",
   286 => x"7f414100",
   287 => x"0800007f",
   288 => x"0603060c",
   289 => x"8000080c",
   290 => x"80808080",
   291 => x"00008080",
   292 => x"07030000",
   293 => x"00000004",
   294 => x"54547420",
   295 => x"0000787c",
   296 => x"44447f7f",
   297 => x"0000387c",
   298 => x"44447c38",
   299 => x"00000044",
   300 => x"44447c38",
   301 => x"00007f7f",
   302 => x"54547c38",
   303 => x"0000185c",
   304 => x"057f7e04",
   305 => x"00000005",
   306 => x"a4a4bc18",
   307 => x"00007cfc",
   308 => x"04047f7f",
   309 => x"0000787c",
   310 => x"7d3d0000",
   311 => x"00000040",
   312 => x"fd808080",
   313 => x"0000007d",
   314 => x"38107f7f",
   315 => x"0000446c",
   316 => x"7f3f0000",
   317 => x"7c000040",
   318 => x"0c180c7c",
   319 => x"0000787c",
   320 => x"04047c7c",
   321 => x"0000787c",
   322 => x"44447c38",
   323 => x"0000387c",
   324 => x"2424fcfc",
   325 => x"0000183c",
   326 => x"24243c18",
   327 => x"0000fcfc",
   328 => x"04047c7c",
   329 => x"0000080c",
   330 => x"54545c48",
   331 => x"00002074",
   332 => x"447f3f04",
   333 => x"00000044",
   334 => x"40407c3c",
   335 => x"00007c7c",
   336 => x"60603c1c",
   337 => x"3c001c3c",
   338 => x"6030607c",
   339 => x"44003c7c",
   340 => x"3810386c",
   341 => x"0000446c",
   342 => x"60e0bc1c",
   343 => x"00001c3c",
   344 => x"5c746444",
   345 => x"0000444c",
   346 => x"773e0808",
   347 => x"00004141",
   348 => x"7f7f0000",
   349 => x"00000000",
   350 => x"3e774141",
   351 => x"02000808",
   352 => x"02030101",
   353 => x"7f000102",
   354 => x"7f7f7f7f",
   355 => x"08007f7f",
   356 => x"3e1c1c08",
   357 => x"7f7f7f3e",
   358 => x"1c3e3e7f",
   359 => x"0008081c",
   360 => x"7c7c1810",
   361 => x"00001018",
   362 => x"7c7c3010",
   363 => x"10001030",
   364 => x"78606030",
   365 => x"4200061e",
   366 => x"3c183c66",
   367 => x"78004266",
   368 => x"c6c26a38",
   369 => x"6000386c",
   370 => x"00600000",
   371 => x"0e006000",
   372 => x"5d5c5b5e",
   373 => x"4c711e0e",
   374 => x"bfdde4c3",
   375 => x"c04bc04d",
   376 => x"02ab741e",
   377 => x"a6c487c7",
   378 => x"c578c048",
   379 => x"48a6c487",
   380 => x"66c478c1",
   381 => x"ee49731e",
   382 => x"86c887df",
   383 => x"ef49e0c0",
   384 => x"a5c487ef",
   385 => x"f0496a4a",
   386 => x"c6f187f0",
   387 => x"c185cb87",
   388 => x"abb7c883",
   389 => x"87c7ff04",
   390 => x"264d2626",
   391 => x"264b264c",
   392 => x"4a711e4f",
   393 => x"5ae1e4c3",
   394 => x"48e1e4c3",
   395 => x"fe4978c7",
   396 => x"4f2687dd",
   397 => x"711e731e",
   398 => x"aab7c04a",
   399 => x"c287d303",
   400 => x"05bfd7e6",
   401 => x"4bc187c4",
   402 => x"4bc087c2",
   403 => x"5bdbe6c2",
   404 => x"e6c287c4",
   405 => x"e6c25adb",
   406 => x"c14abfd7",
   407 => x"a2c0c19a",
   408 => x"87e8ec49",
   409 => x"e6c248fc",
   410 => x"fe78bfd7",
   411 => x"711e87ef",
   412 => x"1e66c44a",
   413 => x"dfff4972",
   414 => x"262687dd",
   415 => x"e6c21e4f",
   416 => x"ff49bfd7",
   417 => x"c387cddc",
   418 => x"e848d5e4",
   419 => x"e4c378bf",
   420 => x"bfec48d1",
   421 => x"d5e4c378",
   422 => x"c3494abf",
   423 => x"b7c899ff",
   424 => x"7148722a",
   425 => x"dde4c3b0",
   426 => x"0e4f2658",
   427 => x"5d5c5b5e",
   428 => x"ff4b710e",
   429 => x"e4c387c7",
   430 => x"50c048d0",
   431 => x"dbff4973",
   432 => x"497087f2",
   433 => x"cb9cc24c",
   434 => x"d2cb49ee",
   435 => x"4d497087",
   436 => x"97d0e4c3",
   437 => x"e4c105bf",
   438 => x"4966d087",
   439 => x"bfd9e4c3",
   440 => x"87d70599",
   441 => x"c34966d4",
   442 => x"99bfd1e4",
   443 => x"7387cc05",
   444 => x"ffdaff49",
   445 => x"02987087",
   446 => x"c187c2c1",
   447 => x"87fdfd4c",
   448 => x"e6ca4975",
   449 => x"02987087",
   450 => x"e4c387c6",
   451 => x"50c148d0",
   452 => x"97d0e4c3",
   453 => x"e4c005bf",
   454 => x"d9e4c387",
   455 => x"66d049bf",
   456 => x"d6ff0599",
   457 => x"d1e4c387",
   458 => x"66d449bf",
   459 => x"caff0599",
   460 => x"ff497387",
   461 => x"7087fdd9",
   462 => x"fefe0598",
   463 => x"fb487487",
   464 => x"5e0e87d7",
   465 => x"0e5d5c5b",
   466 => x"4dc086f4",
   467 => x"7ebfec4c",
   468 => x"c348a6c4",
   469 => x"78bfdde4",
   470 => x"1ec01ec1",
   471 => x"cafd49c7",
   472 => x"7086c887",
   473 => x"87ce0298",
   474 => x"c7fb49ff",
   475 => x"49dac187",
   476 => x"87c0d9ff",
   477 => x"e4c34dc1",
   478 => x"02bf97d0",
   479 => x"f2c087c4",
   480 => x"e4c387d1",
   481 => x"c24bbfd5",
   482 => x"05bfd7e6",
   483 => x"c387ebc0",
   484 => x"d8ff49fd",
   485 => x"fac387de",
   486 => x"d7d8ff49",
   487 => x"c3497387",
   488 => x"1e7199ff",
   489 => x"c5fb49c0",
   490 => x"c8497387",
   491 => x"1e7129b7",
   492 => x"f9fa49c1",
   493 => x"c686c887",
   494 => x"e4c387c3",
   495 => x"9b4bbfd9",
   496 => x"c287dd02",
   497 => x"49bfd3e6",
   498 => x"7087e0c7",
   499 => x"87c40598",
   500 => x"87d24bc0",
   501 => x"c749e0c2",
   502 => x"e6c287c5",
   503 => x"87c658d7",
   504 => x"48d3e6c2",
   505 => x"497378c0",
   506 => x"ce0599c2",
   507 => x"49ebc387",
   508 => x"87c0d7ff",
   509 => x"99c24970",
   510 => x"fb87c202",
   511 => x"c149734c",
   512 => x"87cf0599",
   513 => x"ff49f4c3",
   514 => x"7087e9d6",
   515 => x"0299c249",
   516 => x"fa87c2c0",
   517 => x"c849734c",
   518 => x"87ce0599",
   519 => x"ff49f5c3",
   520 => x"7087d1d6",
   521 => x"0299c249",
   522 => x"e4c387d6",
   523 => x"c002bfe1",
   524 => x"c14887ca",
   525 => x"e5e4c388",
   526 => x"87c2c058",
   527 => x"4dc14cff",
   528 => x"99c44973",
   529 => x"c387ce05",
   530 => x"d5ff49f2",
   531 => x"497087e6",
   532 => x"dc0299c2",
   533 => x"e1e4c387",
   534 => x"c7487ebf",
   535 => x"c003a8b7",
   536 => x"486e87cb",
   537 => x"e4c380c1",
   538 => x"c2c058e5",
   539 => x"c14cfe87",
   540 => x"49fdc34d",
   541 => x"87fcd4ff",
   542 => x"99c24970",
   543 => x"87d5c002",
   544 => x"bfe1e4c3",
   545 => x"87c9c002",
   546 => x"48e1e4c3",
   547 => x"c2c078c0",
   548 => x"c14cfd87",
   549 => x"49fac34d",
   550 => x"87d8d4ff",
   551 => x"99c24970",
   552 => x"87d9c002",
   553 => x"bfe1e4c3",
   554 => x"a8b7c748",
   555 => x"87c9c003",
   556 => x"48e1e4c3",
   557 => x"c2c078c7",
   558 => x"c14cfc87",
   559 => x"acb7c04d",
   560 => x"87d1c003",
   561 => x"c14a66c4",
   562 => x"026a82d8",
   563 => x"6a87c6c0",
   564 => x"7349744b",
   565 => x"c31ec00f",
   566 => x"dac11ef0",
   567 => x"87cbf749",
   568 => x"987086c8",
   569 => x"87e2c002",
   570 => x"c348a6c8",
   571 => x"78bfe1e4",
   572 => x"cb4966c8",
   573 => x"4866c491",
   574 => x"7e708071",
   575 => x"c002bf6e",
   576 => x"bf6e87c8",
   577 => x"4966c84b",
   578 => x"9d750f73",
   579 => x"87c8c002",
   580 => x"bfe1e4c3",
   581 => x"87f7f249",
   582 => x"bfdbe6c2",
   583 => x"87ddc002",
   584 => x"87c7c249",
   585 => x"c0029870",
   586 => x"e4c387d3",
   587 => x"f249bfe1",
   588 => x"49c087dd",
   589 => x"c287fdf3",
   590 => x"c048dbe6",
   591 => x"f38ef478",
   592 => x"5e0e87d7",
   593 => x"0e5d5c5b",
   594 => x"c34c711e",
   595 => x"49bfdde4",
   596 => x"4da1cdc1",
   597 => x"6981d1c1",
   598 => x"029c747e",
   599 => x"a5c487cf",
   600 => x"c37b744b",
   601 => x"49bfdde4",
   602 => x"6e87f6f2",
   603 => x"059c747b",
   604 => x"4bc087c4",
   605 => x"4bc187c2",
   606 => x"f7f24973",
   607 => x"0266d487",
   608 => x"da4987c7",
   609 => x"c24a7087",
   610 => x"c24ac087",
   611 => x"265adfe6",
   612 => x"0087c6f2",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"1e000000",
   616 => x"c8ff4a71",
   617 => x"a17249bf",
   618 => x"1e4f2648",
   619 => x"89bfc8ff",
   620 => x"c0c0c0fe",
   621 => x"01a9c0c0",
   622 => x"4ac087c4",
   623 => x"4ac187c2",
   624 => x"4f264872",
   625 => x"4ad4ff1e",
   626 => x"c848d0ff",
   627 => x"f0c378c5",
   628 => x"c07a717a",
   629 => x"7a7a7a7a",
   630 => x"4f2678c4",
   631 => x"4ad4ff1e",
   632 => x"c848d0ff",
   633 => x"7ac078c5",
   634 => x"7ac0496a",
   635 => x"7a7a7a7a",
   636 => x"487178c4",
   637 => x"5e0e4f26",
   638 => x"0e5d5c5b",
   639 => x"a6cc86e4",
   640 => x"66ecc059",
   641 => x"58a6dc48",
   642 => x"e4c04d70",
   643 => x"e5e4c395",
   644 => x"7ea5d485",
   645 => x"d848a6c4",
   646 => x"66c478a5",
   647 => x"bf6e4cbf",
   648 => x"6d85dc94",
   649 => x"4b66c894",
   650 => x"c0c84ac0",
   651 => x"d4dafd49",
   652 => x"4866c887",
   653 => x"789fc0c1",
   654 => x"c24966c8",
   655 => x"9fbf6e81",
   656 => x"4966c879",
   657 => x"66c481c6",
   658 => x"c8799fbf",
   659 => x"81cc4966",
   660 => x"c8799f6d",
   661 => x"80d44866",
   662 => x"c258a6d0",
   663 => x"cc48ecec",
   664 => x"a1d44966",
   665 => x"7141204a",
   666 => x"87f905aa",
   667 => x"c04866c8",
   668 => x"a6d480ee",
   669 => x"c1edc258",
   670 => x"4966d048",
   671 => x"204aa1c8",
   672 => x"05aa7141",
   673 => x"66c887f9",
   674 => x"80f6c048",
   675 => x"c258a6d8",
   676 => x"d448caed",
   677 => x"e8c04966",
   678 => x"41204aa1",
   679 => x"f905aa71",
   680 => x"4a66d887",
   681 => x"d482f1c0",
   682 => x"81cb4966",
   683 => x"66c85172",
   684 => x"81dec149",
   685 => x"9fd0c0c8",
   686 => x"4966c879",
   687 => x"c881e2c1",
   688 => x"c8799fc0",
   689 => x"eac14966",
   690 => x"799fc181",
   691 => x"c14966c8",
   692 => x"bf6e81ec",
   693 => x"66c8799f",
   694 => x"81eec149",
   695 => x"9fbf66c4",
   696 => x"4966c879",
   697 => x"6d81f0c1",
   698 => x"4b74799f",
   699 => x"9bffffcf",
   700 => x"66c84a73",
   701 => x"81f2c149",
   702 => x"74799f72",
   703 => x"cf2ad04a",
   704 => x"729affff",
   705 => x"4966c84c",
   706 => x"7481f4c1",
   707 => x"c873799f",
   708 => x"f8c14966",
   709 => x"799f7381",
   710 => x"4966c872",
   711 => x"7281fac1",
   712 => x"8ee4799f",
   713 => x"4c264d26",
   714 => x"4f264b26",
   715 => x"53544d69",
   716 => x"6e694d69",
   717 => x"67484d69",
   718 => x"64666172",
   719 => x"6520696c",
   720 => x"30312e00",
   721 => x"20202030",
   722 => x"44650020",
   723 => x"53544d69",
   724 => x"79206966",
   725 => x"20202020",
   726 => x"20202020",
   727 => x"20202020",
   728 => x"20202020",
   729 => x"20202020",
   730 => x"20202020",
   731 => x"20202020",
   732 => x"1e002020",
   733 => x"4b711e73",
   734 => x"d40266d4",
   735 => x"4966c887",
   736 => x"4a7331d8",
   737 => x"a17232c8",
   738 => x"8166cc49",
   739 => x"e1c04871",
   740 => x"4966d087",
   741 => x"c391e4c0",
   742 => x"d881e5e4",
   743 => x"4a6a4aa1",
   744 => x"66c89273",
   745 => x"6981dc82",
   746 => x"cc917249",
   747 => x"89c18166",
   748 => x"f3fd4871",
   749 => x"4a711e87",
   750 => x"ff49d4ff",
   751 => x"c5c848d0",
   752 => x"79d0c278",
   753 => x"797979c0",
   754 => x"79797979",
   755 => x"c0797279",
   756 => x"7966c479",
   757 => x"66c879c0",
   758 => x"cc79c079",
   759 => x"79c07966",
   760 => x"c07966d0",
   761 => x"7966d479",
   762 => x"4f2678c4",
   763 => x"c64a711e",
   764 => x"699749a2",
   765 => x"99f0c349",
   766 => x"1ec01e71",
   767 => x"c01ec11e",
   768 => x"f0fe491e",
   769 => x"49d0c287",
   770 => x"ec87f9f6",
   771 => x"1e4f268e",
   772 => x"1e1e1ec0",
   773 => x"49c11e1e",
   774 => x"c287dafe",
   775 => x"e3f649d0",
   776 => x"268eec87",
   777 => x"4a711e4f",
   778 => x"c848d0ff",
   779 => x"d4ff78c5",
   780 => x"78e0c248",
   781 => x"787878c0",
   782 => x"c0c87878",
   783 => x"fd49721e",
   784 => x"ff87f4d3",
   785 => x"78c448d0",
   786 => x"0e4f2626",
   787 => x"5d5c5b5e",
   788 => x"7186f80e",
   789 => x"4ba2c24a",
   790 => x"c37b97c1",
   791 => x"97c14ca2",
   792 => x"c049a27c",
   793 => x"4da2c451",
   794 => x"c57d97c0",
   795 => x"486e7ea2",
   796 => x"a6c450c0",
   797 => x"78a2c648",
   798 => x"c04866c4",
   799 => x"1e66d850",
   800 => x"49ced2c3",
   801 => x"c887eff5",
   802 => x"49bf9766",
   803 => x"9766c81e",
   804 => x"151e49bf",
   805 => x"49141e49",
   806 => x"1e49131e",
   807 => x"d4fc49c0",
   808 => x"f449c887",
   809 => x"d2c387de",
   810 => x"f8fd49ce",
   811 => x"49d0c287",
   812 => x"e087d1f4",
   813 => x"87ecf98e",
   814 => x"c64a711e",
   815 => x"699749a2",
   816 => x"a2c51e49",
   817 => x"49699749",
   818 => x"49a2c41e",
   819 => x"1e496997",
   820 => x"9749a2c3",
   821 => x"c21e4969",
   822 => x"699749a2",
   823 => x"49c01e49",
   824 => x"c287d2fb",
   825 => x"dbf349d0",
   826 => x"268eec87",
   827 => x"1e731e4f",
   828 => x"a2c24a71",
   829 => x"d04b1149",
   830 => x"c806abb7",
   831 => x"49d1c287",
   832 => x"d587c1f3",
   833 => x"4966c887",
   834 => x"c391e4c0",
   835 => x"c081e5e4",
   836 => x"797381e0",
   837 => x"f249d0c2",
   838 => x"cbf887ea",
   839 => x"1e731e87",
   840 => x"a3c64b71",
   841 => x"49699749",
   842 => x"49a3c51e",
   843 => x"1e496997",
   844 => x"9749a3c4",
   845 => x"c31e4969",
   846 => x"699749a3",
   847 => x"a3c21e49",
   848 => x"49699749",
   849 => x"4aa3c11e",
   850 => x"e8f94912",
   851 => x"49d0c287",
   852 => x"ec87f1f1",
   853 => x"87d0f78e",
   854 => x"5c5b5e0e",
   855 => x"711e0e5d",
   856 => x"c2496e7e",
   857 => x"7997c181",
   858 => x"83c34b6e",
   859 => x"6e7b97c1",
   860 => x"c082c14a",
   861 => x"4c6e7a97",
   862 => x"97c084c4",
   863 => x"c54d6e7c",
   864 => x"6e55c085",
   865 => x"9785c64d",
   866 => x"c01e4d6d",
   867 => x"4c6c971e",
   868 => x"4b6b971e",
   869 => x"4969971e",
   870 => x"f849121e",
   871 => x"d0c287d7",
   872 => x"87e0f049",
   873 => x"fbf58ee8",
   874 => x"5b5e0e87",
   875 => x"ff0e5d5c",
   876 => x"4b7186dc",
   877 => x"1149a3c3",
   878 => x"58a6d448",
   879 => x"c54aa3c4",
   880 => x"699749a3",
   881 => x"9731c849",
   882 => x"71484a6a",
   883 => x"58a6d8b0",
   884 => x"6e7ea3c6",
   885 => x"4d49bf97",
   886 => x"48719dcf",
   887 => x"dc98c0c1",
   888 => x"ec4858a6",
   889 => x"78a3c280",
   890 => x"bf9766c4",
   891 => x"c3059c4c",
   892 => x"4cc0c487",
   893 => x"c01e66d8",
   894 => x"d81e66f8",
   895 => x"1e751e66",
   896 => x"4966e4c0",
   897 => x"d087ecf5",
   898 => x"c0497086",
   899 => x"7459a6e0",
   900 => x"fbc5029c",
   901 => x"66f8c087",
   902 => x"d087c502",
   903 => x"87c55ca6",
   904 => x"c148a6cc",
   905 => x"4b66cc78",
   906 => x"0266f8c0",
   907 => x"f4c087de",
   908 => x"e4c04966",
   909 => x"e5e4c391",
   910 => x"81e0c081",
   911 => x"6948a6c8",
   912 => x"4866cc78",
   913 => x"a8b766c8",
   914 => x"4b87c106",
   915 => x"0566fcc0",
   916 => x"49c887d9",
   917 => x"ee87eded",
   918 => x"497087c2",
   919 => x"ca0599c4",
   920 => x"87f8ed87",
   921 => x"99c44970",
   922 => x"7387f602",
   923 => x"d088c148",
   924 => x"4a7058a6",
   925 => x"c1029b73",
   926 => x"acc187d3",
   927 => x"87c1c102",
   928 => x"4966f4c0",
   929 => x"c391e4c0",
   930 => x"7148e5e4",
   931 => x"58a6cc80",
   932 => x"dc4966c8",
   933 => x"4866d081",
   934 => x"dc05a869",
   935 => x"48a6d087",
   936 => x"c88578c1",
   937 => x"81d84966",
   938 => x"d405ad69",
   939 => x"d44dc087",
   940 => x"80c14866",
   941 => x"c858a6d8",
   942 => x"4866d087",
   943 => x"a6d480c1",
   944 => x"728cc158",
   945 => x"718ac149",
   946 => x"edfe0599",
   947 => x"0266d887",
   948 => x"497387da",
   949 => x"718166dc",
   950 => x"9affc34a",
   951 => x"715aa6d4",
   952 => x"2ab7c84a",
   953 => x"d85aa6d8",
   954 => x"4d7129b7",
   955 => x"49bf976e",
   956 => x"7599f0c3",
   957 => x"d81e71b1",
   958 => x"b7c84966",
   959 => x"dc1e7129",
   960 => x"66dc1e66",
   961 => x"9766d41e",
   962 => x"c01e49bf",
   963 => x"87e5f249",
   964 => x"fcc086d4",
   965 => x"f1c10566",
   966 => x"ea49d087",
   967 => x"f4c087e6",
   968 => x"e4c04966",
   969 => x"e5e4c391",
   970 => x"cc807148",
   971 => x"66c858a6",
   972 => x"6981c849",
   973 => x"87cdc102",
   974 => x"c94966dc",
   975 => x"cc1e7131",
   976 => x"ecfd4966",
   977 => x"86c487ce",
   978 => x"48a6e0c0",
   979 => x"737866cc",
   980 => x"f5c0029b",
   981 => x"cc1ec087",
   982 => x"e9fd4966",
   983 => x"1ec187d8",
   984 => x"fd4966d0",
   985 => x"c887f5e7",
   986 => x"4866dc86",
   987 => x"e0c080c1",
   988 => x"e0c058a6",
   989 => x"c1484966",
   990 => x"a6e4c088",
   991 => x"05997158",
   992 => x"c587d2ff",
   993 => x"e849c987",
   994 => x"9c7487fa",
   995 => x"87c5fa05",
   996 => x"0266fcc0",
   997 => x"d0c287c8",
   998 => x"87e8e849",
   999 => x"c0c287c6",
  1000 => x"87e0e849",
  1001 => x"ed8edcff",
  1002 => x"5e0e87fa",
  1003 => x"0e5d5c5b",
  1004 => x"4c7186e0",
  1005 => x"1149a4c3",
  1006 => x"58a6d448",
  1007 => x"c54aa4c4",
  1008 => x"699749a4",
  1009 => x"9731c849",
  1010 => x"71484a6a",
  1011 => x"58a6d8b0",
  1012 => x"6e7ea4c6",
  1013 => x"4d49bf97",
  1014 => x"48719dcf",
  1015 => x"dc98c0c1",
  1016 => x"ec4858a6",
  1017 => x"78a4c280",
  1018 => x"bf9766c4",
  1019 => x"1e66d84b",
  1020 => x"1e66f4c0",
  1021 => x"751e66d8",
  1022 => x"66e4c01e",
  1023 => x"87f3ed49",
  1024 => x"497086d0",
  1025 => x"59a6e0c0",
  1026 => x"c3059b73",
  1027 => x"4bc0c487",
  1028 => x"efe649c4",
  1029 => x"4966dc87",
  1030 => x"1e7131c9",
  1031 => x"4966f4c0",
  1032 => x"c391e4c0",
  1033 => x"7148e5e4",
  1034 => x"58a6d480",
  1035 => x"fd4966d0",
  1036 => x"c487e1e8",
  1037 => x"029b7386",
  1038 => x"c087ddc4",
  1039 => x"c40266f4",
  1040 => x"c24a7387",
  1041 => x"724ac187",
  1042 => x"66f4c04c",
  1043 => x"cc87d302",
  1044 => x"e0c04966",
  1045 => x"48a6c881",
  1046 => x"66c87869",
  1047 => x"c106aab7",
  1048 => x"9c744c87",
  1049 => x"87d3c202",
  1050 => x"7087f1e5",
  1051 => x"0599c849",
  1052 => x"e7e587ca",
  1053 => x"c8497087",
  1054 => x"87f60299",
  1055 => x"c848d0ff",
  1056 => x"d4ff78c5",
  1057 => x"78f0c248",
  1058 => x"787878c0",
  1059 => x"c0c87878",
  1060 => x"ced2c31e",
  1061 => x"c5c3fd49",
  1062 => x"48d0ff87",
  1063 => x"d2c378c4",
  1064 => x"66d41ece",
  1065 => x"dce5fd49",
  1066 => x"d81ec187",
  1067 => x"e2fd4966",
  1068 => x"86cc87ea",
  1069 => x"c14866dc",
  1070 => x"a6e0c080",
  1071 => x"02abc158",
  1072 => x"cc87f1c0",
  1073 => x"81dc4966",
  1074 => x"694866d0",
  1075 => x"87dc05a8",
  1076 => x"c148a6d0",
  1077 => x"66cc8578",
  1078 => x"6981d849",
  1079 => x"87d405ad",
  1080 => x"66d44dc0",
  1081 => x"d880c148",
  1082 => x"87c858a6",
  1083 => x"c14866d0",
  1084 => x"58a6d480",
  1085 => x"058c8bc1",
  1086 => x"d887edfd",
  1087 => x"87da0266",
  1088 => x"c34966dc",
  1089 => x"a6d499ff",
  1090 => x"4966dc59",
  1091 => x"d829b7c8",
  1092 => x"66dc59a6",
  1093 => x"29b7d849",
  1094 => x"976e4d71",
  1095 => x"f0c349bf",
  1096 => x"71b17599",
  1097 => x"4966d81e",
  1098 => x"7129b7c8",
  1099 => x"1e66dc1e",
  1100 => x"d41e66dc",
  1101 => x"49bf9766",
  1102 => x"e949c01e",
  1103 => x"86d487f7",
  1104 => x"c7029b73",
  1105 => x"e149d087",
  1106 => x"87c687fa",
  1107 => x"e149d0c2",
  1108 => x"9b7387f2",
  1109 => x"87e3fb05",
  1110 => x"c7e78ee0",
  1111 => x"5b5e0e87",
  1112 => x"e40e5d5c",
  1113 => x"cc4a7186",
  1114 => x"ffc048a6",
  1115 => x"c180c478",
  1116 => x"80c478ff",
  1117 => x"c478ffc3",
  1118 => x"c878c080",
  1119 => x"496949a2",
  1120 => x"4d7129c9",
  1121 => x"ebc2029d",
  1122 => x"cc4cc087",
  1123 => x"026b4ba6",
  1124 => x"7487cac2",
  1125 => x"7391c449",
  1126 => x"7e6949a1",
  1127 => x"c448a6c8",
  1128 => x"4966c878",
  1129 => x"1e71916e",
  1130 => x"09751e72",
  1131 => x"d5fdfc4a",
  1132 => x"264a2687",
  1133 => x"58a6c849",
  1134 => x"c0c0c0c4",
  1135 => x"cb01adb7",
  1136 => x"b7ffcf87",
  1137 => x"fdc006a8",
  1138 => x"87ebc087",
  1139 => x"c34866c4",
  1140 => x"a8b7ffff",
  1141 => x"87eec004",
  1142 => x"c74866c4",
  1143 => x"a8b7ffff",
  1144 => x"c887c903",
  1145 => x"b7c54866",
  1146 => x"87da03a8",
  1147 => x"cf4866c4",
  1148 => x"a8b7ffff",
  1149 => x"c887cf06",
  1150 => x"80c14866",
  1151 => x"d058a6cc",
  1152 => x"fe06a8b7",
  1153 => x"66c887db",
  1154 => x"a8b7d048",
  1155 => x"c187ce06",
  1156 => x"c4497484",
  1157 => x"49a17391",
  1158 => x"f6fd0569",
  1159 => x"49a2d487",
  1160 => x"d87966c4",
  1161 => x"66c849a2",
  1162 => x"49a2dc79",
  1163 => x"e0c0796e",
  1164 => x"79c149a2",
  1165 => x"ebe38ee4",
  1166 => x"49c01e87",
  1167 => x"bfede4c3",
  1168 => x"c187c202",
  1169 => x"d1e5c349",
  1170 => x"87c202bf",
  1171 => x"d0ffb1c2",
  1172 => x"78c5c848",
  1173 => x"c348d4ff",
  1174 => x"787178fa",
  1175 => x"c448d0ff",
  1176 => x"1e4f2678",
  1177 => x"4a711e73",
  1178 => x"4966cc1e",
  1179 => x"c391e4c0",
  1180 => x"714be5e4",
  1181 => x"fd497383",
  1182 => x"c487e6d9",
  1183 => x"02987086",
  1184 => x"497387c5",
  1185 => x"fe87d6fb",
  1186 => x"dbe287ef",
  1187 => x"5b5e0e87",
  1188 => x"f40e5d5c",
  1189 => x"c3ddff86",
  1190 => x"c4497087",
  1191 => x"ecc50299",
  1192 => x"48d0ff87",
  1193 => x"ff78c5c8",
  1194 => x"c0c248d4",
  1195 => x"7878c078",
  1196 => x"4d787878",
  1197 => x"c048d4ff",
  1198 => x"a54a7678",
  1199 => x"bfd4ff49",
  1200 => x"d4ff7997",
  1201 => x"6878c048",
  1202 => x"c885c151",
  1203 => x"e304adb7",
  1204 => x"48d0ff87",
  1205 => x"97c678c4",
  1206 => x"a6cc4866",
  1207 => x"d04b7058",
  1208 => x"2bb7c49b",
  1209 => x"e4c04973",
  1210 => x"e5e4c391",
  1211 => x"6981c881",
  1212 => x"c287ca05",
  1213 => x"dbff49d1",
  1214 => x"d0c487ca",
  1215 => x"6697c787",
  1216 => x"f0c3494c",
  1217 => x"05a9d099",
  1218 => x"1e7387cc",
  1219 => x"dbe34972",
  1220 => x"c386c487",
  1221 => x"d0c287f7",
  1222 => x"87c805ac",
  1223 => x"eee34972",
  1224 => x"87e9c387",
  1225 => x"05acecc3",
  1226 => x"1ec087ce",
  1227 => x"49721e73",
  1228 => x"c887d8e4",
  1229 => x"87d5c386",
  1230 => x"05acd1c2",
  1231 => x"1e7387cc",
  1232 => x"f3e54972",
  1233 => x"c386c487",
  1234 => x"c6c387c3",
  1235 => x"87cc05ac",
  1236 => x"49721e73",
  1237 => x"c487d6e6",
  1238 => x"87f1c286",
  1239 => x"05ace0c0",
  1240 => x"1ec087cf",
  1241 => x"721e731e",
  1242 => x"87fde849",
  1243 => x"dcc286cc",
  1244 => x"acc4c387",
  1245 => x"c087d005",
  1246 => x"731ec11e",
  1247 => x"e849721e",
  1248 => x"86cc87e7",
  1249 => x"c087c6c2",
  1250 => x"ce05acf0",
  1251 => x"731ec087",
  1252 => x"f049721e",
  1253 => x"86c887d4",
  1254 => x"c387f2c1",
  1255 => x"ce05acc5",
  1256 => x"731ec187",
  1257 => x"f049721e",
  1258 => x"86c887c0",
  1259 => x"c887dec1",
  1260 => x"87cc05ac",
  1261 => x"49721e73",
  1262 => x"c487dde6",
  1263 => x"87cdc186",
  1264 => x"05acc0c1",
  1265 => x"1ec187d0",
  1266 => x"1e731ec0",
  1267 => x"d8e74972",
  1268 => x"c086cc87",
  1269 => x"9c7487f7",
  1270 => x"7387cc05",
  1271 => x"e449721e",
  1272 => x"86c487fb",
  1273 => x"c887e6c0",
  1274 => x"97c91e66",
  1275 => x"cc1e4966",
  1276 => x"1e496697",
  1277 => x"496697cf",
  1278 => x"6697d21e",
  1279 => x"49c41e49",
  1280 => x"87f1deff",
  1281 => x"d1c286d4",
  1282 => x"f7d6ff49",
  1283 => x"ff8ef487",
  1284 => x"1e87d1dc",
  1285 => x"bfe1d1c3",
  1286 => x"c3b9c149",
  1287 => x"ff59e5d1",
  1288 => x"ffc348d4",
  1289 => x"48d0ff78",
  1290 => x"ff78e1c8",
  1291 => x"78c148d4",
  1292 => x"787131c4",
  1293 => x"c048d0ff",
  1294 => x"4f2678e0",
  1295 => x"d5d1c31e",
  1296 => x"c4dfc31e",
  1297 => x"d8d2fd49",
  1298 => x"7086c487",
  1299 => x"87c30298",
  1300 => x"2687c0ff",
  1301 => x"4b35314f",
  1302 => x"20205a48",
  1303 => x"47464320",
  1304 => x"00000000",
  1305 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
