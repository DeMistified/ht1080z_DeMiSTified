
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"48",x"6e",x"87",x"c4"),
     1 => (x"66",x"c8",x"50",x"c0"),
     2 => (x"c3",x"87",x"c7",x"05"),
     3 => (x"c4",x"48",x"e4",x"e3"),
     4 => (x"85",x"c1",x"78",x"a5"),
     5 => (x"04",x"ad",x"b7",x"c4"),
     6 => (x"c4",x"87",x"c0",x"ff"),
     7 => (x"e3",x"c3",x"87",x"dc"),
     8 => (x"c8",x"48",x"bf",x"f0"),
     9 => (x"d1",x"01",x"a8",x"b7"),
    10 => (x"02",x"ac",x"ca",x"87"),
    11 => (x"ac",x"cd",x"87",x"cc"),
    12 => (x"c0",x"87",x"c7",x"02"),
    13 => (x"c0",x"03",x"ac",x"b7"),
    14 => (x"e3",x"c3",x"87",x"f3"),
    15 => (x"c8",x"4b",x"bf",x"f0"),
    16 => (x"d2",x"03",x"ab",x"b7"),
    17 => (x"f4",x"e3",x"c3",x"87"),
    18 => (x"c0",x"81",x"73",x"49"),
    19 => (x"83",x"c1",x"51",x"e0"),
    20 => (x"04",x"ab",x"b7",x"c8"),
    21 => (x"c3",x"87",x"ee",x"ff"),
    22 => (x"c1",x"48",x"fc",x"e3"),
    23 => (x"cf",x"c1",x"50",x"d2"),
    24 => (x"50",x"cd",x"c1",x"50"),
    25 => (x"80",x"e4",x"50",x"c0"),
    26 => (x"cd",x"c3",x"78",x"c3"),
    27 => (x"f0",x"e3",x"c3",x"87"),
    28 => (x"c1",x"48",x"49",x"bf"),
    29 => (x"f4",x"e3",x"c3",x"80"),
    30 => (x"a0",x"c4",x"48",x"58"),
    31 => (x"c2",x"51",x"74",x"81"),
    32 => (x"f0",x"c0",x"87",x"f8"),
    33 => (x"da",x"04",x"ac",x"b7"),
    34 => (x"b7",x"f9",x"c0",x"87"),
    35 => (x"87",x"d3",x"01",x"ac"),
    36 => (x"bf",x"e8",x"e3",x"c3"),
    37 => (x"74",x"91",x"ca",x"49"),
    38 => (x"8a",x"f0",x"c0",x"4a"),
    39 => (x"48",x"e8",x"e3",x"c3"),
    40 => (x"ca",x"78",x"a1",x"72"),
    41 => (x"c6",x"c0",x"02",x"ac"),
    42 => (x"05",x"ac",x"cd",x"87"),
    43 => (x"c3",x"87",x"cb",x"c2"),
    44 => (x"c3",x"48",x"e4",x"e3"),
    45 => (x"87",x"c2",x"c2",x"78"),
    46 => (x"ac",x"b7",x"f0",x"c0"),
    47 => (x"c0",x"87",x"db",x"04"),
    48 => (x"01",x"ac",x"b7",x"f9"),
    49 => (x"c3",x"87",x"d3",x"c0"),
    50 => (x"49",x"bf",x"ec",x"e3"),
    51 => (x"4a",x"74",x"91",x"d0"),
    52 => (x"c3",x"8a",x"f0",x"c0"),
    53 => (x"72",x"48",x"ec",x"e3"),
    54 => (x"c1",x"c1",x"78",x"a1"),
    55 => (x"c0",x"04",x"ac",x"b7"),
    56 => (x"c6",x"c1",x"87",x"db"),
    57 => (x"c0",x"01",x"ac",x"b7"),
    58 => (x"e3",x"c3",x"87",x"d3"),
    59 => (x"d0",x"49",x"bf",x"ec"),
    60 => (x"c0",x"4a",x"74",x"91"),
    61 => (x"e3",x"c3",x"8a",x"f7"),
    62 => (x"a1",x"72",x"48",x"ec"),
    63 => (x"02",x"ac",x"ca",x"78"),
    64 => (x"cd",x"87",x"c6",x"c0"),
    65 => (x"f1",x"c0",x"05",x"ac"),
    66 => (x"e4",x"e3",x"c3",x"87"),
    67 => (x"c0",x"78",x"c3",x"48"),
    68 => (x"e2",x"c0",x"87",x"e8"),
    69 => (x"c9",x"c0",x"05",x"ac"),
    70 => (x"48",x"a6",x"c4",x"87"),
    71 => (x"c0",x"78",x"fb",x"c0"),
    72 => (x"ac",x"ca",x"87",x"d8"),
    73 => (x"87",x"c6",x"c0",x"02"),
    74 => (x"c0",x"05",x"ac",x"cd"),
    75 => (x"e3",x"c3",x"87",x"c9"),
    76 => (x"78",x"c3",x"48",x"e4"),
    77 => (x"c8",x"87",x"c3",x"c0"),
    78 => (x"b7",x"c0",x"5c",x"a6"),
    79 => (x"c4",x"c0",x"03",x"ac"),
    80 => (x"ca",x"c0",x"48",x"87"),
    81 => (x"02",x"66",x"c4",x"87"),
    82 => (x"48",x"87",x"c6",x"f9"),
    83 => (x"f4",x"99",x"ff",x"c3"),
    84 => (x"87",x"cf",x"f8",x"8e"),
    85 => (x"46",x"4e",x"4f",x"43"),
    86 => (x"4f",x"4d",x"00",x"3d"),
    87 => (x"41",x"4e",x"00",x"44"),
    88 => (x"44",x"00",x"45",x"4d"),
    89 => (x"55",x"41",x"46",x"45"),
    90 => (x"30",x"3d",x"54",x"4c"),
    91 => (x"00",x"21",x"54",x"00"),
    92 => (x"00",x"21",x"5a",x"00"),
    93 => (x"00",x"21",x"5e",x"00"),
    94 => (x"00",x"21",x"63",x"00"),
    95 => (x"d0",x"ff",x"1e",x"00"),
    96 => (x"78",x"c9",x"c8",x"48"),
    97 => (x"d4",x"ff",x"48",x"71"),
    98 => (x"4f",x"26",x"78",x"08"),
    99 => (x"49",x"4a",x"71",x"1e"),
   100 => (x"d0",x"ff",x"87",x"eb"),
   101 => (x"26",x"78",x"c8",x"48"),
   102 => (x"1e",x"73",x"1e",x"4f"),
   103 => (x"e4",x"c3",x"4b",x"71"),
   104 => (x"c3",x"02",x"bf",x"cc"),
   105 => (x"87",x"eb",x"c2",x"87"),
   106 => (x"c8",x"48",x"d0",x"ff"),
   107 => (x"49",x"73",x"78",x"c9"),
   108 => (x"ff",x"b1",x"e0",x"c0"),
   109 => (x"78",x"71",x"48",x"d4"),
   110 => (x"48",x"c0",x"e4",x"c3"),
   111 => (x"66",x"c8",x"78",x"c0"),
   112 => (x"c3",x"87",x"c5",x"02"),
   113 => (x"87",x"c2",x"49",x"ff"),
   114 => (x"e4",x"c3",x"49",x"c0"),
   115 => (x"66",x"cc",x"59",x"c8"),
   116 => (x"c5",x"87",x"c6",x"02"),
   117 => (x"c4",x"4a",x"d5",x"d5"),
   118 => (x"ff",x"ff",x"cf",x"87"),
   119 => (x"cc",x"e4",x"c3",x"4a"),
   120 => (x"cc",x"e4",x"c3",x"5a"),
   121 => (x"c4",x"78",x"c1",x"48"),
   122 => (x"26",x"4d",x"26",x"87"),
   123 => (x"26",x"4b",x"26",x"4c"),
   124 => (x"5b",x"5e",x"0e",x"4f"),
   125 => (x"71",x"0e",x"5d",x"5c"),
   126 => (x"c8",x"e4",x"c3",x"4a"),
   127 => (x"9a",x"72",x"4c",x"bf"),
   128 => (x"49",x"87",x"cb",x"02"),
   129 => (x"c6",x"c2",x"91",x"c8"),
   130 => (x"83",x"71",x"4b",x"cf"),
   131 => (x"ca",x"c2",x"87",x"c4"),
   132 => (x"4d",x"c0",x"4b",x"cf"),
   133 => (x"99",x"74",x"49",x"13"),
   134 => (x"bf",x"c4",x"e4",x"c3"),
   135 => (x"48",x"d4",x"ff",x"b9"),
   136 => (x"b7",x"c1",x"78",x"71"),
   137 => (x"b7",x"c8",x"85",x"2c"),
   138 => (x"87",x"e8",x"04",x"ad"),
   139 => (x"bf",x"c0",x"e4",x"c3"),
   140 => (x"c3",x"80",x"c8",x"48"),
   141 => (x"fe",x"58",x"c4",x"e4"),
   142 => (x"73",x"1e",x"87",x"ef"),
   143 => (x"13",x"4b",x"71",x"1e"),
   144 => (x"cb",x"02",x"9a",x"4a"),
   145 => (x"fe",x"49",x"72",x"87"),
   146 => (x"4a",x"13",x"87",x"e7"),
   147 => (x"87",x"f5",x"05",x"9a"),
   148 => (x"1e",x"87",x"da",x"fe"),
   149 => (x"bf",x"c0",x"e4",x"c3"),
   150 => (x"c0",x"e4",x"c3",x"49"),
   151 => (x"78",x"a1",x"c1",x"48"),
   152 => (x"a9",x"b7",x"c0",x"c4"),
   153 => (x"ff",x"87",x"db",x"03"),
   154 => (x"e4",x"c3",x"48",x"d4"),
   155 => (x"c3",x"78",x"bf",x"c4"),
   156 => (x"49",x"bf",x"c0",x"e4"),
   157 => (x"48",x"c0",x"e4",x"c3"),
   158 => (x"c4",x"78",x"a1",x"c1"),
   159 => (x"04",x"a9",x"b7",x"c0"),
   160 => (x"d0",x"ff",x"87",x"e5"),
   161 => (x"c3",x"78",x"c8",x"48"),
   162 => (x"c0",x"48",x"cc",x"e4"),
   163 => (x"00",x"4f",x"26",x"78"),
   164 => (x"00",x"00",x"00",x"00"),
   165 => (x"00",x"00",x"00",x"00"),
   166 => (x"5f",x"5f",x"00",x"00"),
   167 => (x"00",x"00",x"00",x"00"),
   168 => (x"03",x"00",x"03",x"03"),
   169 => (x"14",x"00",x"00",x"03"),
   170 => (x"7f",x"14",x"7f",x"7f"),
   171 => (x"00",x"00",x"14",x"7f"),
   172 => (x"6b",x"6b",x"2e",x"24"),
   173 => (x"4c",x"00",x"12",x"3a"),
   174 => (x"6c",x"18",x"36",x"6a"),
   175 => (x"30",x"00",x"32",x"56"),
   176 => (x"77",x"59",x"4f",x"7e"),
   177 => (x"00",x"40",x"68",x"3a"),
   178 => (x"03",x"07",x"04",x"00"),
   179 => (x"00",x"00",x"00",x"00"),
   180 => (x"63",x"3e",x"1c",x"00"),
   181 => (x"00",x"00",x"00",x"41"),
   182 => (x"3e",x"63",x"41",x"00"),
   183 => (x"08",x"00",x"00",x"1c"),
   184 => (x"1c",x"1c",x"3e",x"2a"),
   185 => (x"00",x"08",x"2a",x"3e"),
   186 => (x"3e",x"3e",x"08",x"08"),
   187 => (x"00",x"00",x"08",x"08"),
   188 => (x"60",x"e0",x"80",x"00"),
   189 => (x"00",x"00",x"00",x"00"),
   190 => (x"08",x"08",x"08",x"08"),
   191 => (x"00",x"00",x"08",x"08"),
   192 => (x"60",x"60",x"00",x"00"),
   193 => (x"40",x"00",x"00",x"00"),
   194 => (x"0c",x"18",x"30",x"60"),
   195 => (x"00",x"01",x"03",x"06"),
   196 => (x"4d",x"59",x"7f",x"3e"),
   197 => (x"00",x"00",x"3e",x"7f"),
   198 => (x"7f",x"7f",x"06",x"04"),
   199 => (x"00",x"00",x"00",x"00"),
   200 => (x"59",x"71",x"63",x"42"),
   201 => (x"00",x"00",x"46",x"4f"),
   202 => (x"49",x"49",x"63",x"22"),
   203 => (x"18",x"00",x"36",x"7f"),
   204 => (x"7f",x"13",x"16",x"1c"),
   205 => (x"00",x"00",x"10",x"7f"),
   206 => (x"45",x"45",x"67",x"27"),
   207 => (x"00",x"00",x"39",x"7d"),
   208 => (x"49",x"4b",x"7e",x"3c"),
   209 => (x"00",x"00",x"30",x"79"),
   210 => (x"79",x"71",x"01",x"01"),
   211 => (x"00",x"00",x"07",x"0f"),
   212 => (x"49",x"49",x"7f",x"36"),
   213 => (x"00",x"00",x"36",x"7f"),
   214 => (x"69",x"49",x"4f",x"06"),
   215 => (x"00",x"00",x"1e",x"3f"),
   216 => (x"66",x"66",x"00",x"00"),
   217 => (x"00",x"00",x"00",x"00"),
   218 => (x"66",x"e6",x"80",x"00"),
   219 => (x"00",x"00",x"00",x"00"),
   220 => (x"14",x"14",x"08",x"08"),
   221 => (x"00",x"00",x"22",x"22"),
   222 => (x"14",x"14",x"14",x"14"),
   223 => (x"00",x"00",x"14",x"14"),
   224 => (x"14",x"14",x"22",x"22"),
   225 => (x"00",x"00",x"08",x"08"),
   226 => (x"59",x"51",x"03",x"02"),
   227 => (x"3e",x"00",x"06",x"0f"),
   228 => (x"55",x"5d",x"41",x"7f"),
   229 => (x"00",x"00",x"1e",x"1f"),
   230 => (x"09",x"09",x"7f",x"7e"),
   231 => (x"00",x"00",x"7e",x"7f"),
   232 => (x"49",x"49",x"7f",x"7f"),
   233 => (x"00",x"00",x"36",x"7f"),
   234 => (x"41",x"63",x"3e",x"1c"),
   235 => (x"00",x"00",x"41",x"41"),
   236 => (x"63",x"41",x"7f",x"7f"),
   237 => (x"00",x"00",x"1c",x"3e"),
   238 => (x"49",x"49",x"7f",x"7f"),
   239 => (x"00",x"00",x"41",x"41"),
   240 => (x"09",x"09",x"7f",x"7f"),
   241 => (x"00",x"00",x"01",x"01"),
   242 => (x"49",x"41",x"7f",x"3e"),
   243 => (x"00",x"00",x"7a",x"7b"),
   244 => (x"08",x"08",x"7f",x"7f"),
   245 => (x"00",x"00",x"7f",x"7f"),
   246 => (x"7f",x"7f",x"41",x"00"),
   247 => (x"00",x"00",x"00",x"41"),
   248 => (x"40",x"40",x"60",x"20"),
   249 => (x"7f",x"00",x"3f",x"7f"),
   250 => (x"36",x"1c",x"08",x"7f"),
   251 => (x"00",x"00",x"41",x"63"),
   252 => (x"40",x"40",x"7f",x"7f"),
   253 => (x"7f",x"00",x"40",x"40"),
   254 => (x"06",x"0c",x"06",x"7f"),
   255 => (x"7f",x"00",x"7f",x"7f"),
   256 => (x"18",x"0c",x"06",x"7f"),
   257 => (x"00",x"00",x"7f",x"7f"),
   258 => (x"41",x"41",x"7f",x"3e"),
   259 => (x"00",x"00",x"3e",x"7f"),
   260 => (x"09",x"09",x"7f",x"7f"),
   261 => (x"3e",x"00",x"06",x"0f"),
   262 => (x"7f",x"61",x"41",x"7f"),
   263 => (x"00",x"00",x"40",x"7e"),
   264 => (x"19",x"09",x"7f",x"7f"),
   265 => (x"00",x"00",x"66",x"7f"),
   266 => (x"59",x"4d",x"6f",x"26"),
   267 => (x"00",x"00",x"32",x"7b"),
   268 => (x"7f",x"7f",x"01",x"01"),
   269 => (x"00",x"00",x"01",x"01"),
   270 => (x"40",x"40",x"7f",x"3f"),
   271 => (x"00",x"00",x"3f",x"7f"),
   272 => (x"70",x"70",x"3f",x"0f"),
   273 => (x"7f",x"00",x"0f",x"3f"),
   274 => (x"30",x"18",x"30",x"7f"),
   275 => (x"41",x"00",x"7f",x"7f"),
   276 => (x"1c",x"1c",x"36",x"63"),
   277 => (x"01",x"41",x"63",x"36"),
   278 => (x"7c",x"7c",x"06",x"03"),
   279 => (x"61",x"01",x"03",x"06"),
   280 => (x"47",x"4d",x"59",x"71"),
   281 => (x"00",x"00",x"41",x"43"),
   282 => (x"41",x"7f",x"7f",x"00"),
   283 => (x"01",x"00",x"00",x"41"),
   284 => (x"18",x"0c",x"06",x"03"),
   285 => (x"00",x"40",x"60",x"30"),
   286 => (x"7f",x"41",x"41",x"00"),
   287 => (x"08",x"00",x"00",x"7f"),
   288 => (x"06",x"03",x"06",x"0c"),
   289 => (x"80",x"00",x"08",x"0c"),
   290 => (x"80",x"80",x"80",x"80"),
   291 => (x"00",x"00",x"80",x"80"),
   292 => (x"07",x"03",x"00",x"00"),
   293 => (x"00",x"00",x"00",x"04"),
   294 => (x"54",x"54",x"74",x"20"),
   295 => (x"00",x"00",x"78",x"7c"),
   296 => (x"44",x"44",x"7f",x"7f"),
   297 => (x"00",x"00",x"38",x"7c"),
   298 => (x"44",x"44",x"7c",x"38"),
   299 => (x"00",x"00",x"00",x"44"),
   300 => (x"44",x"44",x"7c",x"38"),
   301 => (x"00",x"00",x"7f",x"7f"),
   302 => (x"54",x"54",x"7c",x"38"),
   303 => (x"00",x"00",x"18",x"5c"),
   304 => (x"05",x"7f",x"7e",x"04"),
   305 => (x"00",x"00",x"00",x"05"),
   306 => (x"a4",x"a4",x"bc",x"18"),
   307 => (x"00",x"00",x"7c",x"fc"),
   308 => (x"04",x"04",x"7f",x"7f"),
   309 => (x"00",x"00",x"78",x"7c"),
   310 => (x"7d",x"3d",x"00",x"00"),
   311 => (x"00",x"00",x"00",x"40"),
   312 => (x"fd",x"80",x"80",x"80"),
   313 => (x"00",x"00",x"00",x"7d"),
   314 => (x"38",x"10",x"7f",x"7f"),
   315 => (x"00",x"00",x"44",x"6c"),
   316 => (x"7f",x"3f",x"00",x"00"),
   317 => (x"7c",x"00",x"00",x"40"),
   318 => (x"0c",x"18",x"0c",x"7c"),
   319 => (x"00",x"00",x"78",x"7c"),
   320 => (x"04",x"04",x"7c",x"7c"),
   321 => (x"00",x"00",x"78",x"7c"),
   322 => (x"44",x"44",x"7c",x"38"),
   323 => (x"00",x"00",x"38",x"7c"),
   324 => (x"24",x"24",x"fc",x"fc"),
   325 => (x"00",x"00",x"18",x"3c"),
   326 => (x"24",x"24",x"3c",x"18"),
   327 => (x"00",x"00",x"fc",x"fc"),
   328 => (x"04",x"04",x"7c",x"7c"),
   329 => (x"00",x"00",x"08",x"0c"),
   330 => (x"54",x"54",x"5c",x"48"),
   331 => (x"00",x"00",x"20",x"74"),
   332 => (x"44",x"7f",x"3f",x"04"),
   333 => (x"00",x"00",x"00",x"44"),
   334 => (x"40",x"40",x"7c",x"3c"),
   335 => (x"00",x"00",x"7c",x"7c"),
   336 => (x"60",x"60",x"3c",x"1c"),
   337 => (x"3c",x"00",x"1c",x"3c"),
   338 => (x"60",x"30",x"60",x"7c"),
   339 => (x"44",x"00",x"3c",x"7c"),
   340 => (x"38",x"10",x"38",x"6c"),
   341 => (x"00",x"00",x"44",x"6c"),
   342 => (x"60",x"e0",x"bc",x"1c"),
   343 => (x"00",x"00",x"1c",x"3c"),
   344 => (x"5c",x"74",x"64",x"44"),
   345 => (x"00",x"00",x"44",x"4c"),
   346 => (x"77",x"3e",x"08",x"08"),
   347 => (x"00",x"00",x"41",x"41"),
   348 => (x"7f",x"7f",x"00",x"00"),
   349 => (x"00",x"00",x"00",x"00"),
   350 => (x"3e",x"77",x"41",x"41"),
   351 => (x"02",x"00",x"08",x"08"),
   352 => (x"02",x"03",x"01",x"01"),
   353 => (x"7f",x"00",x"01",x"02"),
   354 => (x"7f",x"7f",x"7f",x"7f"),
   355 => (x"08",x"00",x"7f",x"7f"),
   356 => (x"3e",x"1c",x"1c",x"08"),
   357 => (x"7f",x"7f",x"7f",x"3e"),
   358 => (x"1c",x"3e",x"3e",x"7f"),
   359 => (x"00",x"08",x"08",x"1c"),
   360 => (x"7c",x"7c",x"18",x"10"),
   361 => (x"00",x"00",x"10",x"18"),
   362 => (x"7c",x"7c",x"30",x"10"),
   363 => (x"10",x"00",x"10",x"30"),
   364 => (x"78",x"60",x"60",x"30"),
   365 => (x"42",x"00",x"06",x"1e"),
   366 => (x"3c",x"18",x"3c",x"66"),
   367 => (x"78",x"00",x"42",x"66"),
   368 => (x"c6",x"c2",x"6a",x"38"),
   369 => (x"60",x"00",x"38",x"6c"),
   370 => (x"00",x"60",x"00",x"00"),
   371 => (x"0e",x"00",x"60",x"00"),
   372 => (x"5d",x"5c",x"5b",x"5e"),
   373 => (x"4c",x"71",x"1e",x"0e"),
   374 => (x"bf",x"dd",x"e4",x"c3"),
   375 => (x"c0",x"4b",x"c0",x"4d"),
   376 => (x"02",x"ab",x"74",x"1e"),
   377 => (x"a6",x"c4",x"87",x"c7"),
   378 => (x"c5",x"78",x"c0",x"48"),
   379 => (x"48",x"a6",x"c4",x"87"),
   380 => (x"66",x"c4",x"78",x"c1"),
   381 => (x"ee",x"49",x"73",x"1e"),
   382 => (x"86",x"c8",x"87",x"df"),
   383 => (x"ef",x"49",x"e0",x"c0"),
   384 => (x"a5",x"c4",x"87",x"ef"),
   385 => (x"f0",x"49",x"6a",x"4a"),
   386 => (x"c6",x"f1",x"87",x"f0"),
   387 => (x"c1",x"85",x"cb",x"87"),
   388 => (x"ab",x"b7",x"c8",x"83"),
   389 => (x"87",x"c7",x"ff",x"04"),
   390 => (x"26",x"4d",x"26",x"26"),
   391 => (x"26",x"4b",x"26",x"4c"),
   392 => (x"4a",x"71",x"1e",x"4f"),
   393 => (x"5a",x"e1",x"e4",x"c3"),
   394 => (x"48",x"e1",x"e4",x"c3"),
   395 => (x"fe",x"49",x"78",x"c7"),
   396 => (x"4f",x"26",x"87",x"dd"),
   397 => (x"71",x"1e",x"73",x"1e"),
   398 => (x"aa",x"b7",x"c0",x"4a"),
   399 => (x"c2",x"87",x"d3",x"03"),
   400 => (x"05",x"bf",x"d7",x"e6"),
   401 => (x"4b",x"c1",x"87",x"c4"),
   402 => (x"4b",x"c0",x"87",x"c2"),
   403 => (x"5b",x"db",x"e6",x"c2"),
   404 => (x"e6",x"c2",x"87",x"c4"),
   405 => (x"e6",x"c2",x"5a",x"db"),
   406 => (x"c1",x"4a",x"bf",x"d7"),
   407 => (x"a2",x"c0",x"c1",x"9a"),
   408 => (x"87",x"e8",x"ec",x"49"),
   409 => (x"e6",x"c2",x"48",x"fc"),
   410 => (x"fe",x"78",x"bf",x"d7"),
   411 => (x"71",x"1e",x"87",x"ef"),
   412 => (x"1e",x"66",x"c4",x"4a"),
   413 => (x"df",x"ff",x"49",x"72"),
   414 => (x"26",x"26",x"87",x"dd"),
   415 => (x"e6",x"c2",x"1e",x"4f"),
   416 => (x"ff",x"49",x"bf",x"d7"),
   417 => (x"c3",x"87",x"cd",x"dc"),
   418 => (x"e8",x"48",x"d5",x"e4"),
   419 => (x"e4",x"c3",x"78",x"bf"),
   420 => (x"bf",x"ec",x"48",x"d1"),
   421 => (x"d5",x"e4",x"c3",x"78"),
   422 => (x"c3",x"49",x"4a",x"bf"),
   423 => (x"b7",x"c8",x"99",x"ff"),
   424 => (x"71",x"48",x"72",x"2a"),
   425 => (x"dd",x"e4",x"c3",x"b0"),
   426 => (x"0e",x"4f",x"26",x"58"),
   427 => (x"5d",x"5c",x"5b",x"5e"),
   428 => (x"ff",x"4b",x"71",x"0e"),
   429 => (x"e4",x"c3",x"87",x"c7"),
   430 => (x"50",x"c0",x"48",x"d0"),
   431 => (x"db",x"ff",x"49",x"73"),
   432 => (x"49",x"70",x"87",x"f2"),
   433 => (x"cb",x"9c",x"c2",x"4c"),
   434 => (x"d2",x"cb",x"49",x"ee"),
   435 => (x"4d",x"49",x"70",x"87"),
   436 => (x"97",x"d0",x"e4",x"c3"),
   437 => (x"e4",x"c1",x"05",x"bf"),
   438 => (x"49",x"66",x"d0",x"87"),
   439 => (x"bf",x"d9",x"e4",x"c3"),
   440 => (x"87",x"d7",x"05",x"99"),
   441 => (x"c3",x"49",x"66",x"d4"),
   442 => (x"99",x"bf",x"d1",x"e4"),
   443 => (x"73",x"87",x"cc",x"05"),
   444 => (x"ff",x"da",x"ff",x"49"),
   445 => (x"02",x"98",x"70",x"87"),
   446 => (x"c1",x"87",x"c2",x"c1"),
   447 => (x"87",x"fd",x"fd",x"4c"),
   448 => (x"e6",x"ca",x"49",x"75"),
   449 => (x"02",x"98",x"70",x"87"),
   450 => (x"e4",x"c3",x"87",x"c6"),
   451 => (x"50",x"c1",x"48",x"d0"),
   452 => (x"97",x"d0",x"e4",x"c3"),
   453 => (x"e4",x"c0",x"05",x"bf"),
   454 => (x"d9",x"e4",x"c3",x"87"),
   455 => (x"66",x"d0",x"49",x"bf"),
   456 => (x"d6",x"ff",x"05",x"99"),
   457 => (x"d1",x"e4",x"c3",x"87"),
   458 => (x"66",x"d4",x"49",x"bf"),
   459 => (x"ca",x"ff",x"05",x"99"),
   460 => (x"ff",x"49",x"73",x"87"),
   461 => (x"70",x"87",x"fd",x"d9"),
   462 => (x"fe",x"fe",x"05",x"98"),
   463 => (x"fb",x"48",x"74",x"87"),
   464 => (x"5e",x"0e",x"87",x"d7"),
   465 => (x"0e",x"5d",x"5c",x"5b"),
   466 => (x"4d",x"c0",x"86",x"f4"),
   467 => (x"7e",x"bf",x"ec",x"4c"),
   468 => (x"c3",x"48",x"a6",x"c4"),
   469 => (x"78",x"bf",x"dd",x"e4"),
   470 => (x"1e",x"c0",x"1e",x"c1"),
   471 => (x"ca",x"fd",x"49",x"c7"),
   472 => (x"70",x"86",x"c8",x"87"),
   473 => (x"87",x"ce",x"02",x"98"),
   474 => (x"c7",x"fb",x"49",x"ff"),
   475 => (x"49",x"da",x"c1",x"87"),
   476 => (x"87",x"c0",x"d9",x"ff"),
   477 => (x"e4",x"c3",x"4d",x"c1"),
   478 => (x"02",x"bf",x"97",x"d0"),
   479 => (x"f2",x"c0",x"87",x"c4"),
   480 => (x"e4",x"c3",x"87",x"d1"),
   481 => (x"c2",x"4b",x"bf",x"d5"),
   482 => (x"05",x"bf",x"d7",x"e6"),
   483 => (x"c3",x"87",x"eb",x"c0"),
   484 => (x"d8",x"ff",x"49",x"fd"),
   485 => (x"fa",x"c3",x"87",x"de"),
   486 => (x"d7",x"d8",x"ff",x"49"),
   487 => (x"c3",x"49",x"73",x"87"),
   488 => (x"1e",x"71",x"99",x"ff"),
   489 => (x"c5",x"fb",x"49",x"c0"),
   490 => (x"c8",x"49",x"73",x"87"),
   491 => (x"1e",x"71",x"29",x"b7"),
   492 => (x"f9",x"fa",x"49",x"c1"),
   493 => (x"c6",x"86",x"c8",x"87"),
   494 => (x"e4",x"c3",x"87",x"c3"),
   495 => (x"9b",x"4b",x"bf",x"d9"),
   496 => (x"c2",x"87",x"dd",x"02"),
   497 => (x"49",x"bf",x"d3",x"e6"),
   498 => (x"70",x"87",x"e0",x"c7"),
   499 => (x"87",x"c4",x"05",x"98"),
   500 => (x"87",x"d2",x"4b",x"c0"),
   501 => (x"c7",x"49",x"e0",x"c2"),
   502 => (x"e6",x"c2",x"87",x"c5"),
   503 => (x"87",x"c6",x"58",x"d7"),
   504 => (x"48",x"d3",x"e6",x"c2"),
   505 => (x"49",x"73",x"78",x"c0"),
   506 => (x"ce",x"05",x"99",x"c2"),
   507 => (x"49",x"eb",x"c3",x"87"),
   508 => (x"87",x"c0",x"d7",x"ff"),
   509 => (x"99",x"c2",x"49",x"70"),
   510 => (x"fb",x"87",x"c2",x"02"),
   511 => (x"c1",x"49",x"73",x"4c"),
   512 => (x"87",x"cf",x"05",x"99"),
   513 => (x"ff",x"49",x"f4",x"c3"),
   514 => (x"70",x"87",x"e9",x"d6"),
   515 => (x"02",x"99",x"c2",x"49"),
   516 => (x"fa",x"87",x"c2",x"c0"),
   517 => (x"c8",x"49",x"73",x"4c"),
   518 => (x"87",x"ce",x"05",x"99"),
   519 => (x"ff",x"49",x"f5",x"c3"),
   520 => (x"70",x"87",x"d1",x"d6"),
   521 => (x"02",x"99",x"c2",x"49"),
   522 => (x"e4",x"c3",x"87",x"d6"),
   523 => (x"c0",x"02",x"bf",x"e1"),
   524 => (x"c1",x"48",x"87",x"ca"),
   525 => (x"e5",x"e4",x"c3",x"88"),
   526 => (x"87",x"c2",x"c0",x"58"),
   527 => (x"4d",x"c1",x"4c",x"ff"),
   528 => (x"99",x"c4",x"49",x"73"),
   529 => (x"c3",x"87",x"ce",x"05"),
   530 => (x"d5",x"ff",x"49",x"f2"),
   531 => (x"49",x"70",x"87",x"e6"),
   532 => (x"dc",x"02",x"99",x"c2"),
   533 => (x"e1",x"e4",x"c3",x"87"),
   534 => (x"c7",x"48",x"7e",x"bf"),
   535 => (x"c0",x"03",x"a8",x"b7"),
   536 => (x"48",x"6e",x"87",x"cb"),
   537 => (x"e4",x"c3",x"80",x"c1"),
   538 => (x"c2",x"c0",x"58",x"e5"),
   539 => (x"c1",x"4c",x"fe",x"87"),
   540 => (x"49",x"fd",x"c3",x"4d"),
   541 => (x"87",x"fc",x"d4",x"ff"),
   542 => (x"99",x"c2",x"49",x"70"),
   543 => (x"87",x"d5",x"c0",x"02"),
   544 => (x"bf",x"e1",x"e4",x"c3"),
   545 => (x"87",x"c9",x"c0",x"02"),
   546 => (x"48",x"e1",x"e4",x"c3"),
   547 => (x"c2",x"c0",x"78",x"c0"),
   548 => (x"c1",x"4c",x"fd",x"87"),
   549 => (x"49",x"fa",x"c3",x"4d"),
   550 => (x"87",x"d8",x"d4",x"ff"),
   551 => (x"99",x"c2",x"49",x"70"),
   552 => (x"87",x"d9",x"c0",x"02"),
   553 => (x"bf",x"e1",x"e4",x"c3"),
   554 => (x"a8",x"b7",x"c7",x"48"),
   555 => (x"87",x"c9",x"c0",x"03"),
   556 => (x"48",x"e1",x"e4",x"c3"),
   557 => (x"c2",x"c0",x"78",x"c7"),
   558 => (x"c1",x"4c",x"fc",x"87"),
   559 => (x"ac",x"b7",x"c0",x"4d"),
   560 => (x"87",x"d1",x"c0",x"03"),
   561 => (x"c1",x"4a",x"66",x"c4"),
   562 => (x"02",x"6a",x"82",x"d8"),
   563 => (x"6a",x"87",x"c6",x"c0"),
   564 => (x"73",x"49",x"74",x"4b"),
   565 => (x"c3",x"1e",x"c0",x"0f"),
   566 => (x"da",x"c1",x"1e",x"f0"),
   567 => (x"87",x"cb",x"f7",x"49"),
   568 => (x"98",x"70",x"86",x"c8"),
   569 => (x"87",x"e2",x"c0",x"02"),
   570 => (x"c3",x"48",x"a6",x"c8"),
   571 => (x"78",x"bf",x"e1",x"e4"),
   572 => (x"cb",x"49",x"66",x"c8"),
   573 => (x"48",x"66",x"c4",x"91"),
   574 => (x"7e",x"70",x"80",x"71"),
   575 => (x"c0",x"02",x"bf",x"6e"),
   576 => (x"bf",x"6e",x"87",x"c8"),
   577 => (x"49",x"66",x"c8",x"4b"),
   578 => (x"9d",x"75",x"0f",x"73"),
   579 => (x"87",x"c8",x"c0",x"02"),
   580 => (x"bf",x"e1",x"e4",x"c3"),
   581 => (x"87",x"f7",x"f2",x"49"),
   582 => (x"bf",x"db",x"e6",x"c2"),
   583 => (x"87",x"dd",x"c0",x"02"),
   584 => (x"87",x"c7",x"c2",x"49"),
   585 => (x"c0",x"02",x"98",x"70"),
   586 => (x"e4",x"c3",x"87",x"d3"),
   587 => (x"f2",x"49",x"bf",x"e1"),
   588 => (x"49",x"c0",x"87",x"dd"),
   589 => (x"c2",x"87",x"fd",x"f3"),
   590 => (x"c0",x"48",x"db",x"e6"),
   591 => (x"f3",x"8e",x"f4",x"78"),
   592 => (x"5e",x"0e",x"87",x"d7"),
   593 => (x"0e",x"5d",x"5c",x"5b"),
   594 => (x"c3",x"4c",x"71",x"1e"),
   595 => (x"49",x"bf",x"dd",x"e4"),
   596 => (x"4d",x"a1",x"cd",x"c1"),
   597 => (x"69",x"81",x"d1",x"c1"),
   598 => (x"02",x"9c",x"74",x"7e"),
   599 => (x"a5",x"c4",x"87",x"cf"),
   600 => (x"c3",x"7b",x"74",x"4b"),
   601 => (x"49",x"bf",x"dd",x"e4"),
   602 => (x"6e",x"87",x"f6",x"f2"),
   603 => (x"05",x"9c",x"74",x"7b"),
   604 => (x"4b",x"c0",x"87",x"c4"),
   605 => (x"4b",x"c1",x"87",x"c2"),
   606 => (x"f7",x"f2",x"49",x"73"),
   607 => (x"02",x"66",x"d4",x"87"),
   608 => (x"da",x"49",x"87",x"c7"),
   609 => (x"c2",x"4a",x"70",x"87"),
   610 => (x"c2",x"4a",x"c0",x"87"),
   611 => (x"26",x"5a",x"df",x"e6"),
   612 => (x"00",x"87",x"c6",x"f2"),
   613 => (x"00",x"00",x"00",x"00"),
   614 => (x"00",x"00",x"00",x"00"),
   615 => (x"1e",x"00",x"00",x"00"),
   616 => (x"c8",x"ff",x"4a",x"71"),
   617 => (x"a1",x"72",x"49",x"bf"),
   618 => (x"1e",x"4f",x"26",x"48"),
   619 => (x"89",x"bf",x"c8",x"ff"),
   620 => (x"c0",x"c0",x"c0",x"fe"),
   621 => (x"01",x"a9",x"c0",x"c0"),
   622 => (x"4a",x"c0",x"87",x"c4"),
   623 => (x"4a",x"c1",x"87",x"c2"),
   624 => (x"4f",x"26",x"48",x"72"),
   625 => (x"4a",x"d4",x"ff",x"1e"),
   626 => (x"c8",x"48",x"d0",x"ff"),
   627 => (x"f0",x"c3",x"78",x"c5"),
   628 => (x"c0",x"7a",x"71",x"7a"),
   629 => (x"7a",x"7a",x"7a",x"7a"),
   630 => (x"4f",x"26",x"78",x"c4"),
   631 => (x"4a",x"d4",x"ff",x"1e"),
   632 => (x"c8",x"48",x"d0",x"ff"),
   633 => (x"7a",x"c0",x"78",x"c5"),
   634 => (x"7a",x"c0",x"49",x"6a"),
   635 => (x"7a",x"7a",x"7a",x"7a"),
   636 => (x"48",x"71",x"78",x"c4"),
   637 => (x"5e",x"0e",x"4f",x"26"),
   638 => (x"0e",x"5d",x"5c",x"5b"),
   639 => (x"a6",x"cc",x"86",x"e4"),
   640 => (x"66",x"ec",x"c0",x"59"),
   641 => (x"58",x"a6",x"dc",x"48"),
   642 => (x"e4",x"c0",x"4d",x"70"),
   643 => (x"e5",x"e4",x"c3",x"95"),
   644 => (x"7e",x"a5",x"d4",x"85"),
   645 => (x"d8",x"48",x"a6",x"c4"),
   646 => (x"66",x"c4",x"78",x"a5"),
   647 => (x"bf",x"6e",x"4c",x"bf"),
   648 => (x"6d",x"85",x"dc",x"94"),
   649 => (x"4b",x"66",x"c8",x"94"),
   650 => (x"c0",x"c8",x"4a",x"c0"),
   651 => (x"d4",x"da",x"fd",x"49"),
   652 => (x"48",x"66",x"c8",x"87"),
   653 => (x"78",x"9f",x"c0",x"c1"),
   654 => (x"c2",x"49",x"66",x"c8"),
   655 => (x"9f",x"bf",x"6e",x"81"),
   656 => (x"49",x"66",x"c8",x"79"),
   657 => (x"66",x"c4",x"81",x"c6"),
   658 => (x"c8",x"79",x"9f",x"bf"),
   659 => (x"81",x"cc",x"49",x"66"),
   660 => (x"c8",x"79",x"9f",x"6d"),
   661 => (x"80",x"d4",x"48",x"66"),
   662 => (x"c2",x"58",x"a6",x"d0"),
   663 => (x"cc",x"48",x"ec",x"ec"),
   664 => (x"a1",x"d4",x"49",x"66"),
   665 => (x"71",x"41",x"20",x"4a"),
   666 => (x"87",x"f9",x"05",x"aa"),
   667 => (x"c0",x"48",x"66",x"c8"),
   668 => (x"a6",x"d4",x"80",x"ee"),
   669 => (x"c1",x"ed",x"c2",x"58"),
   670 => (x"49",x"66",x"d0",x"48"),
   671 => (x"20",x"4a",x"a1",x"c8"),
   672 => (x"05",x"aa",x"71",x"41"),
   673 => (x"66",x"c8",x"87",x"f9"),
   674 => (x"80",x"f6",x"c0",x"48"),
   675 => (x"c2",x"58",x"a6",x"d8"),
   676 => (x"d4",x"48",x"ca",x"ed"),
   677 => (x"e8",x"c0",x"49",x"66"),
   678 => (x"41",x"20",x"4a",x"a1"),
   679 => (x"f9",x"05",x"aa",x"71"),
   680 => (x"4a",x"66",x"d8",x"87"),
   681 => (x"d4",x"82",x"f1",x"c0"),
   682 => (x"81",x"cb",x"49",x"66"),
   683 => (x"66",x"c8",x"51",x"72"),
   684 => (x"81",x"de",x"c1",x"49"),
   685 => (x"9f",x"d0",x"c0",x"c8"),
   686 => (x"49",x"66",x"c8",x"79"),
   687 => (x"c8",x"81",x"e2",x"c1"),
   688 => (x"c8",x"79",x"9f",x"c0"),
   689 => (x"ea",x"c1",x"49",x"66"),
   690 => (x"79",x"9f",x"c1",x"81"),
   691 => (x"c1",x"49",x"66",x"c8"),
   692 => (x"bf",x"6e",x"81",x"ec"),
   693 => (x"66",x"c8",x"79",x"9f"),
   694 => (x"81",x"ee",x"c1",x"49"),
   695 => (x"9f",x"bf",x"66",x"c4"),
   696 => (x"49",x"66",x"c8",x"79"),
   697 => (x"6d",x"81",x"f0",x"c1"),
   698 => (x"4b",x"74",x"79",x"9f"),
   699 => (x"9b",x"ff",x"ff",x"cf"),
   700 => (x"66",x"c8",x"4a",x"73"),
   701 => (x"81",x"f2",x"c1",x"49"),
   702 => (x"74",x"79",x"9f",x"72"),
   703 => (x"cf",x"2a",x"d0",x"4a"),
   704 => (x"72",x"9a",x"ff",x"ff"),
   705 => (x"49",x"66",x"c8",x"4c"),
   706 => (x"74",x"81",x"f4",x"c1"),
   707 => (x"c8",x"73",x"79",x"9f"),
   708 => (x"f8",x"c1",x"49",x"66"),
   709 => (x"79",x"9f",x"73",x"81"),
   710 => (x"49",x"66",x"c8",x"72"),
   711 => (x"72",x"81",x"fa",x"c1"),
   712 => (x"8e",x"e4",x"79",x"9f"),
   713 => (x"4c",x"26",x"4d",x"26"),
   714 => (x"4f",x"26",x"4b",x"26"),
   715 => (x"53",x"54",x"4d",x"69"),
   716 => (x"6e",x"69",x"4d",x"69"),
   717 => (x"67",x"48",x"4d",x"69"),
   718 => (x"64",x"66",x"61",x"72"),
   719 => (x"65",x"20",x"69",x"6c"),
   720 => (x"30",x"31",x"2e",x"00"),
   721 => (x"20",x"20",x"20",x"30"),
   722 => (x"44",x"65",x"00",x"20"),
   723 => (x"53",x"54",x"4d",x"69"),
   724 => (x"79",x"20",x"69",x"66"),
   725 => (x"20",x"20",x"20",x"20"),
   726 => (x"20",x"20",x"20",x"20"),
   727 => (x"20",x"20",x"20",x"20"),
   728 => (x"20",x"20",x"20",x"20"),
   729 => (x"20",x"20",x"20",x"20"),
   730 => (x"20",x"20",x"20",x"20"),
   731 => (x"20",x"20",x"20",x"20"),
   732 => (x"1e",x"00",x"20",x"20"),
   733 => (x"4b",x"71",x"1e",x"73"),
   734 => (x"d4",x"02",x"66",x"d4"),
   735 => (x"49",x"66",x"c8",x"87"),
   736 => (x"4a",x"73",x"31",x"d8"),
   737 => (x"a1",x"72",x"32",x"c8"),
   738 => (x"81",x"66",x"cc",x"49"),
   739 => (x"e1",x"c0",x"48",x"71"),
   740 => (x"49",x"66",x"d0",x"87"),
   741 => (x"c3",x"91",x"e4",x"c0"),
   742 => (x"d8",x"81",x"e5",x"e4"),
   743 => (x"4a",x"6a",x"4a",x"a1"),
   744 => (x"66",x"c8",x"92",x"73"),
   745 => (x"69",x"81",x"dc",x"82"),
   746 => (x"cc",x"91",x"72",x"49"),
   747 => (x"89",x"c1",x"81",x"66"),
   748 => (x"f3",x"fd",x"48",x"71"),
   749 => (x"4a",x"71",x"1e",x"87"),
   750 => (x"ff",x"49",x"d4",x"ff"),
   751 => (x"c5",x"c8",x"48",x"d0"),
   752 => (x"79",x"d0",x"c2",x"78"),
   753 => (x"79",x"79",x"79",x"c0"),
   754 => (x"79",x"79",x"79",x"79"),
   755 => (x"c0",x"79",x"72",x"79"),
   756 => (x"79",x"66",x"c4",x"79"),
   757 => (x"66",x"c8",x"79",x"c0"),
   758 => (x"cc",x"79",x"c0",x"79"),
   759 => (x"79",x"c0",x"79",x"66"),
   760 => (x"c0",x"79",x"66",x"d0"),
   761 => (x"79",x"66",x"d4",x"79"),
   762 => (x"4f",x"26",x"78",x"c4"),
   763 => (x"c6",x"4a",x"71",x"1e"),
   764 => (x"69",x"97",x"49",x"a2"),
   765 => (x"99",x"f0",x"c3",x"49"),
   766 => (x"1e",x"c0",x"1e",x"71"),
   767 => (x"c0",x"1e",x"c1",x"1e"),
   768 => (x"f0",x"fe",x"49",x"1e"),
   769 => (x"49",x"d0",x"c2",x"87"),
   770 => (x"ec",x"87",x"f9",x"f6"),
   771 => (x"1e",x"4f",x"26",x"8e"),
   772 => (x"1e",x"1e",x"1e",x"c0"),
   773 => (x"49",x"c1",x"1e",x"1e"),
   774 => (x"c2",x"87",x"da",x"fe"),
   775 => (x"e3",x"f6",x"49",x"d0"),
   776 => (x"26",x"8e",x"ec",x"87"),
   777 => (x"4a",x"71",x"1e",x"4f"),
   778 => (x"c8",x"48",x"d0",x"ff"),
   779 => (x"d4",x"ff",x"78",x"c5"),
   780 => (x"78",x"e0",x"c2",x"48"),
   781 => (x"78",x"78",x"78",x"c0"),
   782 => (x"c0",x"c8",x"78",x"78"),
   783 => (x"fd",x"49",x"72",x"1e"),
   784 => (x"ff",x"87",x"f4",x"d3"),
   785 => (x"78",x"c4",x"48",x"d0"),
   786 => (x"0e",x"4f",x"26",x"26"),
   787 => (x"5d",x"5c",x"5b",x"5e"),
   788 => (x"71",x"86",x"f8",x"0e"),
   789 => (x"4b",x"a2",x"c2",x"4a"),
   790 => (x"c3",x"7b",x"97",x"c1"),
   791 => (x"97",x"c1",x"4c",x"a2"),
   792 => (x"c0",x"49",x"a2",x"7c"),
   793 => (x"4d",x"a2",x"c4",x"51"),
   794 => (x"c5",x"7d",x"97",x"c0"),
   795 => (x"48",x"6e",x"7e",x"a2"),
   796 => (x"a6",x"c4",x"50",x"c0"),
   797 => (x"78",x"a2",x"c6",x"48"),
   798 => (x"c0",x"48",x"66",x"c4"),
   799 => (x"1e",x"66",x"d8",x"50"),
   800 => (x"49",x"ce",x"d2",x"c3"),
   801 => (x"c8",x"87",x"ef",x"f5"),
   802 => (x"49",x"bf",x"97",x"66"),
   803 => (x"97",x"66",x"c8",x"1e"),
   804 => (x"15",x"1e",x"49",x"bf"),
   805 => (x"49",x"14",x"1e",x"49"),
   806 => (x"1e",x"49",x"13",x"1e"),
   807 => (x"d4",x"fc",x"49",x"c0"),
   808 => (x"f4",x"49",x"c8",x"87"),
   809 => (x"d2",x"c3",x"87",x"de"),
   810 => (x"f8",x"fd",x"49",x"ce"),
   811 => (x"49",x"d0",x"c2",x"87"),
   812 => (x"e0",x"87",x"d1",x"f4"),
   813 => (x"87",x"ec",x"f9",x"8e"),
   814 => (x"c6",x"4a",x"71",x"1e"),
   815 => (x"69",x"97",x"49",x"a2"),
   816 => (x"a2",x"c5",x"1e",x"49"),
   817 => (x"49",x"69",x"97",x"49"),
   818 => (x"49",x"a2",x"c4",x"1e"),
   819 => (x"1e",x"49",x"69",x"97"),
   820 => (x"97",x"49",x"a2",x"c3"),
   821 => (x"c2",x"1e",x"49",x"69"),
   822 => (x"69",x"97",x"49",x"a2"),
   823 => (x"49",x"c0",x"1e",x"49"),
   824 => (x"c2",x"87",x"d2",x"fb"),
   825 => (x"db",x"f3",x"49",x"d0"),
   826 => (x"26",x"8e",x"ec",x"87"),
   827 => (x"1e",x"73",x"1e",x"4f"),
   828 => (x"a2",x"c2",x"4a",x"71"),
   829 => (x"d0",x"4b",x"11",x"49"),
   830 => (x"c8",x"06",x"ab",x"b7"),
   831 => (x"49",x"d1",x"c2",x"87"),
   832 => (x"d5",x"87",x"c1",x"f3"),
   833 => (x"49",x"66",x"c8",x"87"),
   834 => (x"c3",x"91",x"e4",x"c0"),
   835 => (x"c0",x"81",x"e5",x"e4"),
   836 => (x"79",x"73",x"81",x"e0"),
   837 => (x"f2",x"49",x"d0",x"c2"),
   838 => (x"cb",x"f8",x"87",x"ea"),
   839 => (x"1e",x"73",x"1e",x"87"),
   840 => (x"a3",x"c6",x"4b",x"71"),
   841 => (x"49",x"69",x"97",x"49"),
   842 => (x"49",x"a3",x"c5",x"1e"),
   843 => (x"1e",x"49",x"69",x"97"),
   844 => (x"97",x"49",x"a3",x"c4"),
   845 => (x"c3",x"1e",x"49",x"69"),
   846 => (x"69",x"97",x"49",x"a3"),
   847 => (x"a3",x"c2",x"1e",x"49"),
   848 => (x"49",x"69",x"97",x"49"),
   849 => (x"4a",x"a3",x"c1",x"1e"),
   850 => (x"e8",x"f9",x"49",x"12"),
   851 => (x"49",x"d0",x"c2",x"87"),
   852 => (x"ec",x"87",x"f1",x"f1"),
   853 => (x"87",x"d0",x"f7",x"8e"),
   854 => (x"5c",x"5b",x"5e",x"0e"),
   855 => (x"71",x"1e",x"0e",x"5d"),
   856 => (x"c2",x"49",x"6e",x"7e"),
   857 => (x"79",x"97",x"c1",x"81"),
   858 => (x"83",x"c3",x"4b",x"6e"),
   859 => (x"6e",x"7b",x"97",x"c1"),
   860 => (x"c0",x"82",x"c1",x"4a"),
   861 => (x"4c",x"6e",x"7a",x"97"),
   862 => (x"97",x"c0",x"84",x"c4"),
   863 => (x"c5",x"4d",x"6e",x"7c"),
   864 => (x"6e",x"55",x"c0",x"85"),
   865 => (x"97",x"85",x"c6",x"4d"),
   866 => (x"c0",x"1e",x"4d",x"6d"),
   867 => (x"4c",x"6c",x"97",x"1e"),
   868 => (x"4b",x"6b",x"97",x"1e"),
   869 => (x"49",x"69",x"97",x"1e"),
   870 => (x"f8",x"49",x"12",x"1e"),
   871 => (x"d0",x"c2",x"87",x"d7"),
   872 => (x"87",x"e0",x"f0",x"49"),
   873 => (x"fb",x"f5",x"8e",x"e8"),
   874 => (x"5b",x"5e",x"0e",x"87"),
   875 => (x"ff",x"0e",x"5d",x"5c"),
   876 => (x"4b",x"71",x"86",x"dc"),
   877 => (x"11",x"49",x"a3",x"c3"),
   878 => (x"58",x"a6",x"d4",x"48"),
   879 => (x"c5",x"4a",x"a3",x"c4"),
   880 => (x"69",x"97",x"49",x"a3"),
   881 => (x"97",x"31",x"c8",x"49"),
   882 => (x"71",x"48",x"4a",x"6a"),
   883 => (x"58",x"a6",x"d8",x"b0"),
   884 => (x"6e",x"7e",x"a3",x"c6"),
   885 => (x"4d",x"49",x"bf",x"97"),
   886 => (x"48",x"71",x"9d",x"cf"),
   887 => (x"dc",x"98",x"c0",x"c1"),
   888 => (x"ec",x"48",x"58",x"a6"),
   889 => (x"78",x"a3",x"c2",x"80"),
   890 => (x"bf",x"97",x"66",x"c4"),
   891 => (x"c3",x"05",x"9c",x"4c"),
   892 => (x"4c",x"c0",x"c4",x"87"),
   893 => (x"c0",x"1e",x"66",x"d8"),
   894 => (x"d8",x"1e",x"66",x"f8"),
   895 => (x"1e",x"75",x"1e",x"66"),
   896 => (x"49",x"66",x"e4",x"c0"),
   897 => (x"d0",x"87",x"ec",x"f5"),
   898 => (x"c0",x"49",x"70",x"86"),
   899 => (x"74",x"59",x"a6",x"e0"),
   900 => (x"fb",x"c5",x"02",x"9c"),
   901 => (x"66",x"f8",x"c0",x"87"),
   902 => (x"d0",x"87",x"c5",x"02"),
   903 => (x"87",x"c5",x"5c",x"a6"),
   904 => (x"c1",x"48",x"a6",x"cc"),
   905 => (x"4b",x"66",x"cc",x"78"),
   906 => (x"02",x"66",x"f8",x"c0"),
   907 => (x"f4",x"c0",x"87",x"de"),
   908 => (x"e4",x"c0",x"49",x"66"),
   909 => (x"e5",x"e4",x"c3",x"91"),
   910 => (x"81",x"e0",x"c0",x"81"),
   911 => (x"69",x"48",x"a6",x"c8"),
   912 => (x"48",x"66",x"cc",x"78"),
   913 => (x"a8",x"b7",x"66",x"c8"),
   914 => (x"4b",x"87",x"c1",x"06"),
   915 => (x"05",x"66",x"fc",x"c0"),
   916 => (x"49",x"c8",x"87",x"d9"),
   917 => (x"ee",x"87",x"ed",x"ed"),
   918 => (x"49",x"70",x"87",x"c2"),
   919 => (x"ca",x"05",x"99",x"c4"),
   920 => (x"87",x"f8",x"ed",x"87"),
   921 => (x"99",x"c4",x"49",x"70"),
   922 => (x"73",x"87",x"f6",x"02"),
   923 => (x"d0",x"88",x"c1",x"48"),
   924 => (x"4a",x"70",x"58",x"a6"),
   925 => (x"c1",x"02",x"9b",x"73"),
   926 => (x"ac",x"c1",x"87",x"d3"),
   927 => (x"87",x"c1",x"c1",x"02"),
   928 => (x"49",x"66",x"f4",x"c0"),
   929 => (x"c3",x"91",x"e4",x"c0"),
   930 => (x"71",x"48",x"e5",x"e4"),
   931 => (x"58",x"a6",x"cc",x"80"),
   932 => (x"dc",x"49",x"66",x"c8"),
   933 => (x"48",x"66",x"d0",x"81"),
   934 => (x"dc",x"05",x"a8",x"69"),
   935 => (x"48",x"a6",x"d0",x"87"),
   936 => (x"c8",x"85",x"78",x"c1"),
   937 => (x"81",x"d8",x"49",x"66"),
   938 => (x"d4",x"05",x"ad",x"69"),
   939 => (x"d4",x"4d",x"c0",x"87"),
   940 => (x"80",x"c1",x"48",x"66"),
   941 => (x"c8",x"58",x"a6",x"d8"),
   942 => (x"48",x"66",x"d0",x"87"),
   943 => (x"a6",x"d4",x"80",x"c1"),
   944 => (x"72",x"8c",x"c1",x"58"),
   945 => (x"71",x"8a",x"c1",x"49"),
   946 => (x"ed",x"fe",x"05",x"99"),
   947 => (x"02",x"66",x"d8",x"87"),
   948 => (x"49",x"73",x"87",x"da"),
   949 => (x"71",x"81",x"66",x"dc"),
   950 => (x"9a",x"ff",x"c3",x"4a"),
   951 => (x"71",x"5a",x"a6",x"d4"),
   952 => (x"2a",x"b7",x"c8",x"4a"),
   953 => (x"d8",x"5a",x"a6",x"d8"),
   954 => (x"4d",x"71",x"29",x"b7"),
   955 => (x"49",x"bf",x"97",x"6e"),
   956 => (x"75",x"99",x"f0",x"c3"),
   957 => (x"d8",x"1e",x"71",x"b1"),
   958 => (x"b7",x"c8",x"49",x"66"),
   959 => (x"dc",x"1e",x"71",x"29"),
   960 => (x"66",x"dc",x"1e",x"66"),
   961 => (x"97",x"66",x"d4",x"1e"),
   962 => (x"c0",x"1e",x"49",x"bf"),
   963 => (x"87",x"e5",x"f2",x"49"),
   964 => (x"fc",x"c0",x"86",x"d4"),
   965 => (x"f1",x"c1",x"05",x"66"),
   966 => (x"ea",x"49",x"d0",x"87"),
   967 => (x"f4",x"c0",x"87",x"e6"),
   968 => (x"e4",x"c0",x"49",x"66"),
   969 => (x"e5",x"e4",x"c3",x"91"),
   970 => (x"cc",x"80",x"71",x"48"),
   971 => (x"66",x"c8",x"58",x"a6"),
   972 => (x"69",x"81",x"c8",x"49"),
   973 => (x"87",x"cd",x"c1",x"02"),
   974 => (x"c9",x"49",x"66",x"dc"),
   975 => (x"cc",x"1e",x"71",x"31"),
   976 => (x"ec",x"fd",x"49",x"66"),
   977 => (x"86",x"c4",x"87",x"ce"),
   978 => (x"48",x"a6",x"e0",x"c0"),
   979 => (x"73",x"78",x"66",x"cc"),
   980 => (x"f5",x"c0",x"02",x"9b"),
   981 => (x"cc",x"1e",x"c0",x"87"),
   982 => (x"e9",x"fd",x"49",x"66"),
   983 => (x"1e",x"c1",x"87",x"d8"),
   984 => (x"fd",x"49",x"66",x"d0"),
   985 => (x"c8",x"87",x"f5",x"e7"),
   986 => (x"48",x"66",x"dc",x"86"),
   987 => (x"e0",x"c0",x"80",x"c1"),
   988 => (x"e0",x"c0",x"58",x"a6"),
   989 => (x"c1",x"48",x"49",x"66"),
   990 => (x"a6",x"e4",x"c0",x"88"),
   991 => (x"05",x"99",x"71",x"58"),
   992 => (x"c5",x"87",x"d2",x"ff"),
   993 => (x"e8",x"49",x"c9",x"87"),
   994 => (x"9c",x"74",x"87",x"fa"),
   995 => (x"87",x"c5",x"fa",x"05"),
   996 => (x"02",x"66",x"fc",x"c0"),
   997 => (x"d0",x"c2",x"87",x"c8"),
   998 => (x"87",x"e8",x"e8",x"49"),
   999 => (x"c0",x"c2",x"87",x"c6"),
  1000 => (x"87",x"e0",x"e8",x"49"),
  1001 => (x"ed",x"8e",x"dc",x"ff"),
  1002 => (x"5e",x"0e",x"87",x"fa"),
  1003 => (x"0e",x"5d",x"5c",x"5b"),
  1004 => (x"4c",x"71",x"86",x"e0"),
  1005 => (x"11",x"49",x"a4",x"c3"),
  1006 => (x"58",x"a6",x"d4",x"48"),
  1007 => (x"c5",x"4a",x"a4",x"c4"),
  1008 => (x"69",x"97",x"49",x"a4"),
  1009 => (x"97",x"31",x"c8",x"49"),
  1010 => (x"71",x"48",x"4a",x"6a"),
  1011 => (x"58",x"a6",x"d8",x"b0"),
  1012 => (x"6e",x"7e",x"a4",x"c6"),
  1013 => (x"4d",x"49",x"bf",x"97"),
  1014 => (x"48",x"71",x"9d",x"cf"),
  1015 => (x"dc",x"98",x"c0",x"c1"),
  1016 => (x"ec",x"48",x"58",x"a6"),
  1017 => (x"78",x"a4",x"c2",x"80"),
  1018 => (x"bf",x"97",x"66",x"c4"),
  1019 => (x"1e",x"66",x"d8",x"4b"),
  1020 => (x"1e",x"66",x"f4",x"c0"),
  1021 => (x"75",x"1e",x"66",x"d8"),
  1022 => (x"66",x"e4",x"c0",x"1e"),
  1023 => (x"87",x"f3",x"ed",x"49"),
  1024 => (x"49",x"70",x"86",x"d0"),
  1025 => (x"59",x"a6",x"e0",x"c0"),
  1026 => (x"c3",x"05",x"9b",x"73"),
  1027 => (x"4b",x"c0",x"c4",x"87"),
  1028 => (x"ef",x"e6",x"49",x"c4"),
  1029 => (x"49",x"66",x"dc",x"87"),
  1030 => (x"1e",x"71",x"31",x"c9"),
  1031 => (x"49",x"66",x"f4",x"c0"),
  1032 => (x"c3",x"91",x"e4",x"c0"),
  1033 => (x"71",x"48",x"e5",x"e4"),
  1034 => (x"58",x"a6",x"d4",x"80"),
  1035 => (x"fd",x"49",x"66",x"d0"),
  1036 => (x"c4",x"87",x"e1",x"e8"),
  1037 => (x"02",x"9b",x"73",x"86"),
  1038 => (x"c0",x"87",x"dd",x"c4"),
  1039 => (x"c4",x"02",x"66",x"f4"),
  1040 => (x"c2",x"4a",x"73",x"87"),
  1041 => (x"72",x"4a",x"c1",x"87"),
  1042 => (x"66",x"f4",x"c0",x"4c"),
  1043 => (x"cc",x"87",x"d3",x"02"),
  1044 => (x"e0",x"c0",x"49",x"66"),
  1045 => (x"48",x"a6",x"c8",x"81"),
  1046 => (x"66",x"c8",x"78",x"69"),
  1047 => (x"c1",x"06",x"aa",x"b7"),
  1048 => (x"9c",x"74",x"4c",x"87"),
  1049 => (x"87",x"d3",x"c2",x"02"),
  1050 => (x"70",x"87",x"f1",x"e5"),
  1051 => (x"05",x"99",x"c8",x"49"),
  1052 => (x"e7",x"e5",x"87",x"ca"),
  1053 => (x"c8",x"49",x"70",x"87"),
  1054 => (x"87",x"f6",x"02",x"99"),
  1055 => (x"c8",x"48",x"d0",x"ff"),
  1056 => (x"d4",x"ff",x"78",x"c5"),
  1057 => (x"78",x"f0",x"c2",x"48"),
  1058 => (x"78",x"78",x"78",x"c0"),
  1059 => (x"c0",x"c8",x"78",x"78"),
  1060 => (x"ce",x"d2",x"c3",x"1e"),
  1061 => (x"c5",x"c3",x"fd",x"49"),
  1062 => (x"48",x"d0",x"ff",x"87"),
  1063 => (x"d2",x"c3",x"78",x"c4"),
  1064 => (x"66",x"d4",x"1e",x"ce"),
  1065 => (x"dc",x"e5",x"fd",x"49"),
  1066 => (x"d8",x"1e",x"c1",x"87"),
  1067 => (x"e2",x"fd",x"49",x"66"),
  1068 => (x"86",x"cc",x"87",x"ea"),
  1069 => (x"c1",x"48",x"66",x"dc"),
  1070 => (x"a6",x"e0",x"c0",x"80"),
  1071 => (x"02",x"ab",x"c1",x"58"),
  1072 => (x"cc",x"87",x"f1",x"c0"),
  1073 => (x"81",x"dc",x"49",x"66"),
  1074 => (x"69",x"48",x"66",x"d0"),
  1075 => (x"87",x"dc",x"05",x"a8"),
  1076 => (x"c1",x"48",x"a6",x"d0"),
  1077 => (x"66",x"cc",x"85",x"78"),
  1078 => (x"69",x"81",x"d8",x"49"),
  1079 => (x"87",x"d4",x"05",x"ad"),
  1080 => (x"66",x"d4",x"4d",x"c0"),
  1081 => (x"d8",x"80",x"c1",x"48"),
  1082 => (x"87",x"c8",x"58",x"a6"),
  1083 => (x"c1",x"48",x"66",x"d0"),
  1084 => (x"58",x"a6",x"d4",x"80"),
  1085 => (x"05",x"8c",x"8b",x"c1"),
  1086 => (x"d8",x"87",x"ed",x"fd"),
  1087 => (x"87",x"da",x"02",x"66"),
  1088 => (x"c3",x"49",x"66",x"dc"),
  1089 => (x"a6",x"d4",x"99",x"ff"),
  1090 => (x"49",x"66",x"dc",x"59"),
  1091 => (x"d8",x"29",x"b7",x"c8"),
  1092 => (x"66",x"dc",x"59",x"a6"),
  1093 => (x"29",x"b7",x"d8",x"49"),
  1094 => (x"97",x"6e",x"4d",x"71"),
  1095 => (x"f0",x"c3",x"49",x"bf"),
  1096 => (x"71",x"b1",x"75",x"99"),
  1097 => (x"49",x"66",x"d8",x"1e"),
  1098 => (x"71",x"29",x"b7",x"c8"),
  1099 => (x"1e",x"66",x"dc",x"1e"),
  1100 => (x"d4",x"1e",x"66",x"dc"),
  1101 => (x"49",x"bf",x"97",x"66"),
  1102 => (x"e9",x"49",x"c0",x"1e"),
  1103 => (x"86",x"d4",x"87",x"f7"),
  1104 => (x"c7",x"02",x"9b",x"73"),
  1105 => (x"e1",x"49",x"d0",x"87"),
  1106 => (x"87",x"c6",x"87",x"fa"),
  1107 => (x"e1",x"49",x"d0",x"c2"),
  1108 => (x"9b",x"73",x"87",x"f2"),
  1109 => (x"87",x"e3",x"fb",x"05"),
  1110 => (x"c7",x"e7",x"8e",x"e0"),
  1111 => (x"5b",x"5e",x"0e",x"87"),
  1112 => (x"e4",x"0e",x"5d",x"5c"),
  1113 => (x"cc",x"4a",x"71",x"86"),
  1114 => (x"ff",x"c0",x"48",x"a6"),
  1115 => (x"c1",x"80",x"c4",x"78"),
  1116 => (x"80",x"c4",x"78",x"ff"),
  1117 => (x"c4",x"78",x"ff",x"c3"),
  1118 => (x"c8",x"78",x"c0",x"80"),
  1119 => (x"49",x"69",x"49",x"a2"),
  1120 => (x"4d",x"71",x"29",x"c9"),
  1121 => (x"eb",x"c2",x"02",x"9d"),
  1122 => (x"cc",x"4c",x"c0",x"87"),
  1123 => (x"02",x"6b",x"4b",x"a6"),
  1124 => (x"74",x"87",x"ca",x"c2"),
  1125 => (x"73",x"91",x"c4",x"49"),
  1126 => (x"7e",x"69",x"49",x"a1"),
  1127 => (x"c4",x"48",x"a6",x"c8"),
  1128 => (x"49",x"66",x"c8",x"78"),
  1129 => (x"1e",x"71",x"91",x"6e"),
  1130 => (x"09",x"75",x"1e",x"72"),
  1131 => (x"d5",x"fd",x"fc",x"4a"),
  1132 => (x"26",x"4a",x"26",x"87"),
  1133 => (x"58",x"a6",x"c8",x"49"),
  1134 => (x"c0",x"c0",x"c0",x"c4"),
  1135 => (x"cb",x"01",x"ad",x"b7"),
  1136 => (x"b7",x"ff",x"cf",x"87"),
  1137 => (x"fd",x"c0",x"06",x"a8"),
  1138 => (x"87",x"eb",x"c0",x"87"),
  1139 => (x"c3",x"48",x"66",x"c4"),
  1140 => (x"a8",x"b7",x"ff",x"ff"),
  1141 => (x"87",x"ee",x"c0",x"04"),
  1142 => (x"c7",x"48",x"66",x"c4"),
  1143 => (x"a8",x"b7",x"ff",x"ff"),
  1144 => (x"c8",x"87",x"c9",x"03"),
  1145 => (x"b7",x"c5",x"48",x"66"),
  1146 => (x"87",x"da",x"03",x"a8"),
  1147 => (x"cf",x"48",x"66",x"c4"),
  1148 => (x"a8",x"b7",x"ff",x"ff"),
  1149 => (x"c8",x"87",x"cf",x"06"),
  1150 => (x"80",x"c1",x"48",x"66"),
  1151 => (x"d0",x"58",x"a6",x"cc"),
  1152 => (x"fe",x"06",x"a8",x"b7"),
  1153 => (x"66",x"c8",x"87",x"db"),
  1154 => (x"a8",x"b7",x"d0",x"48"),
  1155 => (x"c1",x"87",x"ce",x"06"),
  1156 => (x"c4",x"49",x"74",x"84"),
  1157 => (x"49",x"a1",x"73",x"91"),
  1158 => (x"f6",x"fd",x"05",x"69"),
  1159 => (x"49",x"a2",x"d4",x"87"),
  1160 => (x"d8",x"79",x"66",x"c4"),
  1161 => (x"66",x"c8",x"49",x"a2"),
  1162 => (x"49",x"a2",x"dc",x"79"),
  1163 => (x"e0",x"c0",x"79",x"6e"),
  1164 => (x"79",x"c1",x"49",x"a2"),
  1165 => (x"eb",x"e3",x"8e",x"e4"),
  1166 => (x"49",x"c0",x"1e",x"87"),
  1167 => (x"bf",x"ed",x"e4",x"c3"),
  1168 => (x"c1",x"87",x"c2",x"02"),
  1169 => (x"d1",x"e5",x"c3",x"49"),
  1170 => (x"87",x"c2",x"02",x"bf"),
  1171 => (x"d0",x"ff",x"b1",x"c2"),
  1172 => (x"78",x"c5",x"c8",x"48"),
  1173 => (x"c3",x"48",x"d4",x"ff"),
  1174 => (x"78",x"71",x"78",x"fa"),
  1175 => (x"c4",x"48",x"d0",x"ff"),
  1176 => (x"1e",x"4f",x"26",x"78"),
  1177 => (x"4a",x"71",x"1e",x"73"),
  1178 => (x"49",x"66",x"cc",x"1e"),
  1179 => (x"c3",x"91",x"e4",x"c0"),
  1180 => (x"71",x"4b",x"e5",x"e4"),
  1181 => (x"fd",x"49",x"73",x"83"),
  1182 => (x"c4",x"87",x"e6",x"d9"),
  1183 => (x"02",x"98",x"70",x"86"),
  1184 => (x"49",x"73",x"87",x"c5"),
  1185 => (x"fe",x"87",x"d6",x"fb"),
  1186 => (x"db",x"e2",x"87",x"ef"),
  1187 => (x"5b",x"5e",x"0e",x"87"),
  1188 => (x"f4",x"0e",x"5d",x"5c"),
  1189 => (x"c3",x"dd",x"ff",x"86"),
  1190 => (x"c4",x"49",x"70",x"87"),
  1191 => (x"ec",x"c5",x"02",x"99"),
  1192 => (x"48",x"d0",x"ff",x"87"),
  1193 => (x"ff",x"78",x"c5",x"c8"),
  1194 => (x"c0",x"c2",x"48",x"d4"),
  1195 => (x"78",x"78",x"c0",x"78"),
  1196 => (x"4d",x"78",x"78",x"78"),
  1197 => (x"c0",x"48",x"d4",x"ff"),
  1198 => (x"a5",x"4a",x"76",x"78"),
  1199 => (x"bf",x"d4",x"ff",x"49"),
  1200 => (x"d4",x"ff",x"79",x"97"),
  1201 => (x"68",x"78",x"c0",x"48"),
  1202 => (x"c8",x"85",x"c1",x"51"),
  1203 => (x"e3",x"04",x"ad",x"b7"),
  1204 => (x"48",x"d0",x"ff",x"87"),
  1205 => (x"97",x"c6",x"78",x"c4"),
  1206 => (x"a6",x"cc",x"48",x"66"),
  1207 => (x"d0",x"4b",x"70",x"58"),
  1208 => (x"2b",x"b7",x"c4",x"9b"),
  1209 => (x"e4",x"c0",x"49",x"73"),
  1210 => (x"e5",x"e4",x"c3",x"91"),
  1211 => (x"69",x"81",x"c8",x"81"),
  1212 => (x"c2",x"87",x"ca",x"05"),
  1213 => (x"db",x"ff",x"49",x"d1"),
  1214 => (x"d0",x"c4",x"87",x"ca"),
  1215 => (x"66",x"97",x"c7",x"87"),
  1216 => (x"f0",x"c3",x"49",x"4c"),
  1217 => (x"05",x"a9",x"d0",x"99"),
  1218 => (x"1e",x"73",x"87",x"cc"),
  1219 => (x"db",x"e3",x"49",x"72"),
  1220 => (x"c3",x"86",x"c4",x"87"),
  1221 => (x"d0",x"c2",x"87",x"f7"),
  1222 => (x"87",x"c8",x"05",x"ac"),
  1223 => (x"ee",x"e3",x"49",x"72"),
  1224 => (x"87",x"e9",x"c3",x"87"),
  1225 => (x"05",x"ac",x"ec",x"c3"),
  1226 => (x"1e",x"c0",x"87",x"ce"),
  1227 => (x"49",x"72",x"1e",x"73"),
  1228 => (x"c8",x"87",x"d8",x"e4"),
  1229 => (x"87",x"d5",x"c3",x"86"),
  1230 => (x"05",x"ac",x"d1",x"c2"),
  1231 => (x"1e",x"73",x"87",x"cc"),
  1232 => (x"f3",x"e5",x"49",x"72"),
  1233 => (x"c3",x"86",x"c4",x"87"),
  1234 => (x"c6",x"c3",x"87",x"c3"),
  1235 => (x"87",x"cc",x"05",x"ac"),
  1236 => (x"49",x"72",x"1e",x"73"),
  1237 => (x"c4",x"87",x"d6",x"e6"),
  1238 => (x"87",x"f1",x"c2",x"86"),
  1239 => (x"05",x"ac",x"e0",x"c0"),
  1240 => (x"1e",x"c0",x"87",x"cf"),
  1241 => (x"72",x"1e",x"73",x"1e"),
  1242 => (x"87",x"fd",x"e8",x"49"),
  1243 => (x"dc",x"c2",x"86",x"cc"),
  1244 => (x"ac",x"c4",x"c3",x"87"),
  1245 => (x"c0",x"87",x"d0",x"05"),
  1246 => (x"73",x"1e",x"c1",x"1e"),
  1247 => (x"e8",x"49",x"72",x"1e"),
  1248 => (x"86",x"cc",x"87",x"e7"),
  1249 => (x"c0",x"87",x"c6",x"c2"),
  1250 => (x"ce",x"05",x"ac",x"f0"),
  1251 => (x"73",x"1e",x"c0",x"87"),
  1252 => (x"f0",x"49",x"72",x"1e"),
  1253 => (x"86",x"c8",x"87",x"d4"),
  1254 => (x"c3",x"87",x"f2",x"c1"),
  1255 => (x"ce",x"05",x"ac",x"c5"),
  1256 => (x"73",x"1e",x"c1",x"87"),
  1257 => (x"f0",x"49",x"72",x"1e"),
  1258 => (x"86",x"c8",x"87",x"c0"),
  1259 => (x"c8",x"87",x"de",x"c1"),
  1260 => (x"87",x"cc",x"05",x"ac"),
  1261 => (x"49",x"72",x"1e",x"73"),
  1262 => (x"c4",x"87",x"dd",x"e6"),
  1263 => (x"87",x"cd",x"c1",x"86"),
  1264 => (x"05",x"ac",x"c0",x"c1"),
  1265 => (x"1e",x"c1",x"87",x"d0"),
  1266 => (x"1e",x"73",x"1e",x"c0"),
  1267 => (x"d8",x"e7",x"49",x"72"),
  1268 => (x"c0",x"86",x"cc",x"87"),
  1269 => (x"9c",x"74",x"87",x"f7"),
  1270 => (x"73",x"87",x"cc",x"05"),
  1271 => (x"e4",x"49",x"72",x"1e"),
  1272 => (x"86",x"c4",x"87",x"fb"),
  1273 => (x"c8",x"87",x"e6",x"c0"),
  1274 => (x"97",x"c9",x"1e",x"66"),
  1275 => (x"cc",x"1e",x"49",x"66"),
  1276 => (x"1e",x"49",x"66",x"97"),
  1277 => (x"49",x"66",x"97",x"cf"),
  1278 => (x"66",x"97",x"d2",x"1e"),
  1279 => (x"49",x"c4",x"1e",x"49"),
  1280 => (x"87",x"f1",x"de",x"ff"),
  1281 => (x"d1",x"c2",x"86",x"d4"),
  1282 => (x"f7",x"d6",x"ff",x"49"),
  1283 => (x"ff",x"8e",x"f4",x"87"),
  1284 => (x"1e",x"87",x"d1",x"dc"),
  1285 => (x"bf",x"e1",x"d1",x"c3"),
  1286 => (x"c3",x"b9",x"c1",x"49"),
  1287 => (x"ff",x"59",x"e5",x"d1"),
  1288 => (x"ff",x"c3",x"48",x"d4"),
  1289 => (x"48",x"d0",x"ff",x"78"),
  1290 => (x"ff",x"78",x"e1",x"c8"),
  1291 => (x"78",x"c1",x"48",x"d4"),
  1292 => (x"78",x"71",x"31",x"c4"),
  1293 => (x"c0",x"48",x"d0",x"ff"),
  1294 => (x"4f",x"26",x"78",x"e0"),
  1295 => (x"d5",x"d1",x"c3",x"1e"),
  1296 => (x"c4",x"df",x"c3",x"1e"),
  1297 => (x"d8",x"d2",x"fd",x"49"),
  1298 => (x"70",x"86",x"c4",x"87"),
  1299 => (x"87",x"c3",x"02",x"98"),
  1300 => (x"26",x"87",x"c0",x"ff"),
  1301 => (x"4b",x"35",x"31",x"4f"),
  1302 => (x"20",x"20",x"5a",x"48"),
  1303 => (x"47",x"46",x"43",x"20"),
  1304 => (x"00",x"00",x"00",x"00"),
  1305 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

