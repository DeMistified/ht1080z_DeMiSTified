library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f0e5c387",
    12 => x"86c0c64e",
    13 => x"49f0e5c3",
    14 => x"48e8d1c3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c0eb",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"731e4f26",
    53 => x"029a721e",
    54 => x"c087e7c0",
    55 => x"724bc148",
    56 => x"87d106a9",
    57 => x"c9068272",
    58 => x"72837387",
    59 => x"87f401a9",
    60 => x"b2c187c3",
    61 => x"03a9723a",
    62 => x"07807389",
    63 => x"052b2ac1",
    64 => x"4b2687f3",
    65 => x"751e4f26",
    66 => x"714dc41e",
    67 => x"ff04a1b7",
    68 => x"c381c1b9",
    69 => x"b77207bd",
    70 => x"baff04a2",
    71 => x"bdc182c1",
    72 => x"87eefe07",
    73 => x"ff042dc1",
    74 => x"0780c1b8",
    75 => x"b9ff042d",
    76 => x"260781c1",
    77 => x"1e4f264d",
    78 => x"66c44a71",
    79 => x"88c14849",
    80 => x"7158a6c8",
    81 => x"87d40299",
    82 => x"d4ff4812",
    83 => x"66c47808",
    84 => x"88c14849",
    85 => x"7158a6c8",
    86 => x"87ec0599",
    87 => x"711e4f26",
    88 => x"4966c44a",
    89 => x"c888c148",
    90 => x"997158a6",
    91 => x"ff87d602",
    92 => x"ffc348d4",
    93 => x"c4526878",
    94 => x"c1484966",
    95 => x"58a6c888",
    96 => x"ea059971",
    97 => x"1e4f2687",
    98 => x"d4ff1e73",
    99 => x"7bffc34b",
   100 => x"ffc34a6b",
   101 => x"c8496b7b",
   102 => x"c3b17232",
   103 => x"4a6b7bff",
   104 => x"b27131c8",
   105 => x"6b7bffc3",
   106 => x"7232c849",
   107 => x"c44871b1",
   108 => x"264d2687",
   109 => x"264b264c",
   110 => x"5b5e0e4f",
   111 => x"710e5d5c",
   112 => x"4cd4ff4a",
   113 => x"ffc34972",
   114 => x"c37c7199",
   115 => x"05bfe8d1",
   116 => x"66d087c8",
   117 => x"d430c948",
   118 => x"66d058a6",
   119 => x"c329d849",
   120 => x"7c7199ff",
   121 => x"d04966d0",
   122 => x"99ffc329",
   123 => x"66d07c71",
   124 => x"c329c849",
   125 => x"7c7199ff",
   126 => x"c34966d0",
   127 => x"7c7199ff",
   128 => x"29d04972",
   129 => x"7199ffc3",
   130 => x"c94b6c7c",
   131 => x"c34dfff0",
   132 => x"d005abff",
   133 => x"7cffc387",
   134 => x"8dc14b6c",
   135 => x"c387c602",
   136 => x"f002abff",
   137 => x"fe487387",
   138 => x"c01e87c7",
   139 => x"48d4ff49",
   140 => x"c178ffc3",
   141 => x"b7c8c381",
   142 => x"87f104a9",
   143 => x"731e4f26",
   144 => x"c487e71e",
   145 => x"c04bdff8",
   146 => x"f0ffc01e",
   147 => x"fd49f7c1",
   148 => x"86c487e7",
   149 => x"c005a8c1",
   150 => x"d4ff87ea",
   151 => x"78ffc348",
   152 => x"c0c0c0c1",
   153 => x"c01ec0c0",
   154 => x"e9c1f0e1",
   155 => x"87c9fd49",
   156 => x"987086c4",
   157 => x"ff87ca05",
   158 => x"ffc348d4",
   159 => x"cb48c178",
   160 => x"87e6fe87",
   161 => x"fe058bc1",
   162 => x"48c087fd",
   163 => x"1e87e6fc",
   164 => x"d4ff1e73",
   165 => x"78ffc348",
   166 => x"1ec04bd3",
   167 => x"c1f0ffc0",
   168 => x"d4fc49c1",
   169 => x"7086c487",
   170 => x"87ca0598",
   171 => x"c348d4ff",
   172 => x"48c178ff",
   173 => x"f1fd87cb",
   174 => x"058bc187",
   175 => x"c087dbff",
   176 => x"87f1fb48",
   177 => x"5c5b5e0e",
   178 => x"4cd4ff0e",
   179 => x"c687dbfd",
   180 => x"e1c01eea",
   181 => x"49c8c1f0",
   182 => x"c487defb",
   183 => x"02a8c186",
   184 => x"eafe87c8",
   185 => x"c148c087",
   186 => x"dafa87e2",
   187 => x"cf497087",
   188 => x"c699ffff",
   189 => x"c802a9ea",
   190 => x"87d3fe87",
   191 => x"cbc148c0",
   192 => x"7cffc387",
   193 => x"fc4bf1c0",
   194 => x"987087f4",
   195 => x"87ebc002",
   196 => x"ffc01ec0",
   197 => x"49fac1f0",
   198 => x"c487defa",
   199 => x"05987086",
   200 => x"ffc387d9",
   201 => x"c3496c7c",
   202 => x"7c7c7cff",
   203 => x"99c0c17c",
   204 => x"c187c402",
   205 => x"c087d548",
   206 => x"c287d148",
   207 => x"87c405ab",
   208 => x"87c848c0",
   209 => x"fe058bc1",
   210 => x"48c087fd",
   211 => x"1e87e4f9",
   212 => x"d1c31e73",
   213 => x"78c148e8",
   214 => x"d0ff4bc7",
   215 => x"fb78c248",
   216 => x"d0ff87c8",
   217 => x"c078c348",
   218 => x"d0e5c01e",
   219 => x"f949c0c1",
   220 => x"86c487c7",
   221 => x"c105a8c1",
   222 => x"abc24b87",
   223 => x"c087c505",
   224 => x"87f9c048",
   225 => x"ff058bc1",
   226 => x"f7fc87d0",
   227 => x"ecd1c387",
   228 => x"05987058",
   229 => x"1ec187cd",
   230 => x"c1f0ffc0",
   231 => x"d8f849d0",
   232 => x"ff86c487",
   233 => x"ffc348d4",
   234 => x"87dec478",
   235 => x"58f0d1c3",
   236 => x"c248d0ff",
   237 => x"48d4ff78",
   238 => x"c178ffc3",
   239 => x"87f5f748",
   240 => x"5c5b5e0e",
   241 => x"4a710e5d",
   242 => x"ff4dffc3",
   243 => x"7c754cd4",
   244 => x"c448d0ff",
   245 => x"7c7578c3",
   246 => x"ffc01e72",
   247 => x"49d8c1f0",
   248 => x"c487d6f7",
   249 => x"02987086",
   250 => x"48c187c5",
   251 => x"7587f0c0",
   252 => x"7cfec37c",
   253 => x"d41ec0c8",
   254 => x"faf44966",
   255 => x"7586c487",
   256 => x"757c757c",
   257 => x"e0dad87c",
   258 => x"6c7c754b",
   259 => x"c5059949",
   260 => x"058bc187",
   261 => x"7c7587f3",
   262 => x"c248d0ff",
   263 => x"f648c078",
   264 => x"5e0e87cf",
   265 => x"0e5d5c5b",
   266 => x"4cc04b71",
   267 => x"dfcdeec5",
   268 => x"48d4ff4a",
   269 => x"6878ffc3",
   270 => x"a9fec349",
   271 => x"87fdc005",
   272 => x"9b734d70",
   273 => x"d087cc02",
   274 => x"49731e66",
   275 => x"c487cff4",
   276 => x"ff87d686",
   277 => x"d1c448d0",
   278 => x"7dffc378",
   279 => x"c14866d0",
   280 => x"58a6d488",
   281 => x"f0059870",
   282 => x"48d4ff87",
   283 => x"7878ffc3",
   284 => x"c5059b73",
   285 => x"48d0ff87",
   286 => x"4ac178d0",
   287 => x"058ac14c",
   288 => x"7487eefe",
   289 => x"87e9f448",
   290 => x"711e731e",
   291 => x"ff4bc04a",
   292 => x"ffc348d4",
   293 => x"48d0ff78",
   294 => x"ff78c3c4",
   295 => x"ffc348d4",
   296 => x"c01e7278",
   297 => x"d1c1f0ff",
   298 => x"87cdf449",
   299 => x"987086c4",
   300 => x"c887d205",
   301 => x"66cc1ec0",
   302 => x"87e6fd49",
   303 => x"4b7086c4",
   304 => x"c248d0ff",
   305 => x"f3487378",
   306 => x"5e0e87eb",
   307 => x"0e5d5c5b",
   308 => x"ffc01ec0",
   309 => x"49c9c1f0",
   310 => x"d287def3",
   311 => x"f0d1c31e",
   312 => x"87fefc49",
   313 => x"4cc086c8",
   314 => x"b7d284c1",
   315 => x"87f804ac",
   316 => x"97f0d1c3",
   317 => x"c0c349bf",
   318 => x"a9c0c199",
   319 => x"87e7c005",
   320 => x"97f7d1c3",
   321 => x"31d049bf",
   322 => x"97f8d1c3",
   323 => x"32c84abf",
   324 => x"d1c3b172",
   325 => x"4abf97f9",
   326 => x"cf4c71b1",
   327 => x"9cffffff",
   328 => x"34ca84c1",
   329 => x"c387e7c1",
   330 => x"bf97f9d1",
   331 => x"c631c149",
   332 => x"fad1c399",
   333 => x"c74abf97",
   334 => x"b1722ab7",
   335 => x"97f5d1c3",
   336 => x"cf4d4abf",
   337 => x"f6d1c39d",
   338 => x"c34abf97",
   339 => x"c332ca9a",
   340 => x"bf97f7d1",
   341 => x"7333c24b",
   342 => x"f8d1c3b2",
   343 => x"c34bbf97",
   344 => x"b7c69bc0",
   345 => x"c2b2732b",
   346 => x"7148c181",
   347 => x"c1497030",
   348 => x"70307548",
   349 => x"c14c724d",
   350 => x"c8947184",
   351 => x"06adb7c0",
   352 => x"34c187cc",
   353 => x"c0c82db7",
   354 => x"ff01adb7",
   355 => x"487487f4",
   356 => x"0e87def0",
   357 => x"5d5c5b5e",
   358 => x"c386f80e",
   359 => x"c048d6da",
   360 => x"ced2c378",
   361 => x"fb49c01e",
   362 => x"86c487de",
   363 => x"c5059870",
   364 => x"c948c087",
   365 => x"4dc087ce",
   366 => x"fac07ec1",
   367 => x"c349bfe1",
   368 => x"714ac4d3",
   369 => x"e1ea4bc8",
   370 => x"05987087",
   371 => x"7ec087c2",
   372 => x"bfddfac0",
   373 => x"e0d3c349",
   374 => x"4bc8714a",
   375 => x"7087cbea",
   376 => x"87c20598",
   377 => x"026e7ec0",
   378 => x"c387fdc0",
   379 => x"4dbfd4d9",
   380 => x"9fccdac3",
   381 => x"c5487ebf",
   382 => x"05a8ead6",
   383 => x"d9c387c7",
   384 => x"ce4dbfd4",
   385 => x"ca486e87",
   386 => x"02a8d5e9",
   387 => x"48c087c5",
   388 => x"c387f1c7",
   389 => x"751eced2",
   390 => x"87ecf949",
   391 => x"987086c4",
   392 => x"c087c505",
   393 => x"87dcc748",
   394 => x"bfddfac0",
   395 => x"e0d3c349",
   396 => x"4bc8714a",
   397 => x"7087f3e8",
   398 => x"87c80598",
   399 => x"48d6dac3",
   400 => x"87da78c1",
   401 => x"bfe1fac0",
   402 => x"c4d3c349",
   403 => x"4bc8714a",
   404 => x"7087d7e8",
   405 => x"c5c00298",
   406 => x"c648c087",
   407 => x"dac387e6",
   408 => x"49bf97cc",
   409 => x"05a9d5c1",
   410 => x"c387cdc0",
   411 => x"bf97cdda",
   412 => x"a9eac249",
   413 => x"87c5c002",
   414 => x"c7c648c0",
   415 => x"ced2c387",
   416 => x"487ebf97",
   417 => x"02a8e9c3",
   418 => x"6e87cec0",
   419 => x"a8ebc348",
   420 => x"87c5c002",
   421 => x"ebc548c0",
   422 => x"d9d2c387",
   423 => x"9949bf97",
   424 => x"87ccc005",
   425 => x"97dad2c3",
   426 => x"a9c249bf",
   427 => x"87c5c002",
   428 => x"cfc548c0",
   429 => x"dbd2c387",
   430 => x"c348bf97",
   431 => x"7058d2da",
   432 => x"88c1484c",
   433 => x"58d6dac3",
   434 => x"97dcd2c3",
   435 => x"817549bf",
   436 => x"97ddd2c3",
   437 => x"32c84abf",
   438 => x"c37ea172",
   439 => x"6e48e3de",
   440 => x"ded2c378",
   441 => x"c848bf97",
   442 => x"dac358a6",
   443 => x"c202bfd6",
   444 => x"fac087d4",
   445 => x"c349bfdd",
   446 => x"714ae0d3",
   447 => x"e9e54bc8",
   448 => x"02987087",
   449 => x"c087c5c0",
   450 => x"87f8c348",
   451 => x"bfcedac3",
   452 => x"f7dec34c",
   453 => x"f3d2c35c",
   454 => x"c849bf97",
   455 => x"f2d2c331",
   456 => x"a14abf97",
   457 => x"f4d2c349",
   458 => x"d04abf97",
   459 => x"49a17232",
   460 => x"97f5d2c3",
   461 => x"32d84abf",
   462 => x"c449a172",
   463 => x"dec39166",
   464 => x"c381bfe3",
   465 => x"c359ebde",
   466 => x"bf97fbd2",
   467 => x"c332c84a",
   468 => x"bf97fad2",
   469 => x"c34aa24b",
   470 => x"bf97fcd2",
   471 => x"7333d04b",
   472 => x"d2c34aa2",
   473 => x"4bbf97fd",
   474 => x"33d89bcf",
   475 => x"c34aa273",
   476 => x"c35aefde",
   477 => x"4abfebde",
   478 => x"92748ac2",
   479 => x"48efdec3",
   480 => x"c178a172",
   481 => x"d2c387ca",
   482 => x"49bf97e0",
   483 => x"d2c331c8",
   484 => x"4abf97df",
   485 => x"dac349a1",
   486 => x"dac359de",
   487 => x"c549bfda",
   488 => x"81ffc731",
   489 => x"dec329c9",
   490 => x"d2c359f7",
   491 => x"4abf97e5",
   492 => x"d2c332c8",
   493 => x"4bbf97e4",
   494 => x"66c44aa2",
   495 => x"c3826e92",
   496 => x"c35af3de",
   497 => x"c048ebde",
   498 => x"e7dec378",
   499 => x"78a17248",
   500 => x"48f7dec3",
   501 => x"bfebdec3",
   502 => x"fbdec378",
   503 => x"efdec348",
   504 => x"dac378bf",
   505 => x"c002bfd6",
   506 => x"487487c9",
   507 => x"7e7030c4",
   508 => x"c387c9c0",
   509 => x"48bff3de",
   510 => x"7e7030c4",
   511 => x"48dadac3",
   512 => x"48c1786e",
   513 => x"4d268ef8",
   514 => x"4b264c26",
   515 => x"5e0e4f26",
   516 => x"0e5d5c5b",
   517 => x"dac34a71",
   518 => x"cb02bfd6",
   519 => x"c74b7287",
   520 => x"c14c722b",
   521 => x"87c99cff",
   522 => x"2bc84b72",
   523 => x"ffc34c72",
   524 => x"e3dec39c",
   525 => x"fac083bf",
   526 => x"02abbfd9",
   527 => x"fac087d9",
   528 => x"d2c35bdd",
   529 => x"49731ece",
   530 => x"c487fdf0",
   531 => x"05987086",
   532 => x"48c087c5",
   533 => x"c387e6c0",
   534 => x"02bfd6da",
   535 => x"497487d2",
   536 => x"d2c391c4",
   537 => x"4d6981ce",
   538 => x"ffffffcf",
   539 => x"87cb9dff",
   540 => x"91c24974",
   541 => x"81ced2c3",
   542 => x"754d699f",
   543 => x"87c6fe48",
   544 => x"5c5b5e0e",
   545 => x"711e0e5d",
   546 => x"c11ec04d",
   547 => x"87edd049",
   548 => x"4c7086c4",
   549 => x"c2c1029c",
   550 => x"dedac387",
   551 => x"ff49754a",
   552 => x"7087ecde",
   553 => x"f2c00298",
   554 => x"754a7487",
   555 => x"ff4bcb49",
   556 => x"7087d1df",
   557 => x"e2c00298",
   558 => x"741ec087",
   559 => x"87c7029c",
   560 => x"c048a6c4",
   561 => x"c487c578",
   562 => x"78c148a6",
   563 => x"cf4966c4",
   564 => x"86c487eb",
   565 => x"059c4c70",
   566 => x"7487fefe",
   567 => x"e5fc2648",
   568 => x"5b5e0e87",
   569 => x"1e0e5d5c",
   570 => x"059b4b71",
   571 => x"48c087c5",
   572 => x"c887e5c1",
   573 => x"7dc04da3",
   574 => x"c70266d4",
   575 => x"9766d487",
   576 => x"87c505bf",
   577 => x"cfc148c0",
   578 => x"4966d487",
   579 => x"7087f1fd",
   580 => x"c1029c4c",
   581 => x"a4dc87c0",
   582 => x"da7d6949",
   583 => x"a3c449a4",
   584 => x"7a699f4a",
   585 => x"bfd6dac3",
   586 => x"d487d202",
   587 => x"699f49a4",
   588 => x"ffffc049",
   589 => x"d0487199",
   590 => x"c27e7030",
   591 => x"6e7ec087",
   592 => x"806a4849",
   593 => x"7bc07a70",
   594 => x"6a49a3cc",
   595 => x"49a3d079",
   596 => x"48c179c0",
   597 => x"48c087c2",
   598 => x"87eafa26",
   599 => x"5c5b5e0e",
   600 => x"4c710e5d",
   601 => x"cac1029c",
   602 => x"49a4c887",
   603 => x"c2c10269",
   604 => x"4a66d087",
   605 => x"d482496c",
   606 => x"66d05aa6",
   607 => x"dac3b94d",
   608 => x"ff4abfd2",
   609 => x"719972ba",
   610 => x"e4c00299",
   611 => x"4ba4c487",
   612 => x"f9f9496b",
   613 => x"c37b7087",
   614 => x"49bfceda",
   615 => x"7c71816c",
   616 => x"dac3b975",
   617 => x"ff4abfd2",
   618 => x"719972ba",
   619 => x"dcff0599",
   620 => x"f97c7587",
   621 => x"731e87d0",
   622 => x"9b4b711e",
   623 => x"c887c702",
   624 => x"056949a3",
   625 => x"48c087c5",
   626 => x"c387f7c0",
   627 => x"4abfe7de",
   628 => x"6949a3c4",
   629 => x"c389c249",
   630 => x"91bfceda",
   631 => x"c34aa271",
   632 => x"49bfd2da",
   633 => x"a271996b",
   634 => x"ddfac04a",
   635 => x"1e66c85a",
   636 => x"d3ea4972",
   637 => x"7086c487",
   638 => x"87c40598",
   639 => x"87c248c0",
   640 => x"c5f848c1",
   641 => x"1e731e87",
   642 => x"029b4b71",
   643 => x"a3c887c7",
   644 => x"c5056949",
   645 => x"c048c087",
   646 => x"dec387f7",
   647 => x"c44abfe7",
   648 => x"496949a3",
   649 => x"dac389c2",
   650 => x"7191bfce",
   651 => x"dac34aa2",
   652 => x"6b49bfd2",
   653 => x"4aa27199",
   654 => x"5addfac0",
   655 => x"721e66c8",
   656 => x"87fce549",
   657 => x"987086c4",
   658 => x"c087c405",
   659 => x"c187c248",
   660 => x"87f6f648",
   661 => x"5c5b5e0e",
   662 => x"711e0e5d",
   663 => x"4c66d44b",
   664 => x"9b732cc9",
   665 => x"87cfc102",
   666 => x"6949a3c8",
   667 => x"87c7c102",
   668 => x"d44da3d0",
   669 => x"dac37d66",
   670 => x"ff49bfd2",
   671 => x"994a6bb9",
   672 => x"03ac717e",
   673 => x"7bc087cd",
   674 => x"4aa3cc7d",
   675 => x"6a49a3c4",
   676 => x"7287c279",
   677 => x"029c748c",
   678 => x"1e4987dd",
   679 => x"fbfa4973",
   680 => x"d486c487",
   681 => x"ffc74966",
   682 => x"87cb0299",
   683 => x"1eced2c3",
   684 => x"c1fc4973",
   685 => x"2686c487",
   686 => x"0e87cbf5",
   687 => x"5d5c5b5e",
   688 => x"d086f00e",
   689 => x"e4c059a6",
   690 => x"66cc4b66",
   691 => x"4887ca02",
   692 => x"7e7080c8",
   693 => x"c505bf6e",
   694 => x"c348c087",
   695 => x"66cc87ec",
   696 => x"7384d04c",
   697 => x"48a6c449",
   698 => x"66c4786c",
   699 => x"6e80c481",
   700 => x"66c878bf",
   701 => x"87c606a9",
   702 => x"8966c449",
   703 => x"b7c04b71",
   704 => x"87c401ab",
   705 => x"87c2c348",
   706 => x"c74866c4",
   707 => x"7e7098ff",
   708 => x"c9c1026e",
   709 => x"49c0c887",
   710 => x"4a71896e",
   711 => x"4dced2c3",
   712 => x"b773856e",
   713 => x"87c106aa",
   714 => x"4849724a",
   715 => x"708066c4",
   716 => x"498b727c",
   717 => x"99718ac1",
   718 => x"c087d902",
   719 => x"154866e0",
   720 => x"66e0c050",
   721 => x"c080c148",
   722 => x"7258a6e4",
   723 => x"718ac149",
   724 => x"87e70599",
   725 => x"66d01ec1",
   726 => x"87c0f849",
   727 => x"b7c086c4",
   728 => x"e3c106ab",
   729 => x"66e0c087",
   730 => x"b7ffc74d",
   731 => x"e2c006ab",
   732 => x"d01e7587",
   733 => x"fdf84966",
   734 => x"85c0c887",
   735 => x"c0c8486c",
   736 => x"c87c7080",
   737 => x"1ec18bc0",
   738 => x"f74966d4",
   739 => x"86c887ce",
   740 => x"c387eec0",
   741 => x"d01eced2",
   742 => x"d9f84966",
   743 => x"c386c487",
   744 => x"734aced2",
   745 => x"806c4849",
   746 => x"49737c70",
   747 => x"99718bc1",
   748 => x"1287ce02",
   749 => x"85c17d97",
   750 => x"8bc14973",
   751 => x"f2059971",
   752 => x"abb7c087",
   753 => x"87e1fe01",
   754 => x"8ef048c1",
   755 => x"0e87f7f0",
   756 => x"5d5c5b5e",
   757 => x"9b4b710e",
   758 => x"c887c702",
   759 => x"056d4da3",
   760 => x"48ff87c5",
   761 => x"d087fdc0",
   762 => x"496c4ca3",
   763 => x"0599ffc7",
   764 => x"026c87d8",
   765 => x"1ec187c9",
   766 => x"dff54973",
   767 => x"c386c487",
   768 => x"731eced2",
   769 => x"87eef649",
   770 => x"4a6c86c4",
   771 => x"c404aa6d",
   772 => x"cf48ff87",
   773 => x"7ca2c187",
   774 => x"ffc74972",
   775 => x"ced2c399",
   776 => x"48699781",
   777 => x"1e87dfef",
   778 => x"4b711e73",
   779 => x"e4c0029b",
   780 => x"fbdec387",
   781 => x"c24a735b",
   782 => x"cedac38a",
   783 => x"c39249bf",
   784 => x"48bfe7de",
   785 => x"dec38072",
   786 => x"487158ff",
   787 => x"dac330c4",
   788 => x"edc058de",
   789 => x"f7dec387",
   790 => x"ebdec348",
   791 => x"dec378bf",
   792 => x"dec348fb",
   793 => x"c378bfef",
   794 => x"02bfd6da",
   795 => x"dac387c9",
   796 => x"c449bfce",
   797 => x"c387c731",
   798 => x"49bff3de",
   799 => x"dac331c4",
   800 => x"c5ee59de",
   801 => x"5b5e0e87",
   802 => x"4a710e5c",
   803 => x"9a724bc0",
   804 => x"87e1c002",
   805 => x"9f49a2da",
   806 => x"dac34b69",
   807 => x"cf02bfd6",
   808 => x"49a2d487",
   809 => x"4c49699f",
   810 => x"9cffffc0",
   811 => x"87c234d0",
   812 => x"49744cc0",
   813 => x"fd4973b3",
   814 => x"cbed87ed",
   815 => x"5b5e0e87",
   816 => x"f40e5d5c",
   817 => x"c04a7186",
   818 => x"029a727e",
   819 => x"d2c387d8",
   820 => x"78c048ca",
   821 => x"48c2d2c3",
   822 => x"bffbdec3",
   823 => x"c6d2c378",
   824 => x"f7dec348",
   825 => x"dac378bf",
   826 => x"50c048eb",
   827 => x"bfdadac3",
   828 => x"cad2c349",
   829 => x"aa714abf",
   830 => x"87cac403",
   831 => x"99cf4972",
   832 => x"87eac005",
   833 => x"48d9fac0",
   834 => x"bfc2d2c3",
   835 => x"ced2c378",
   836 => x"c2d2c31e",
   837 => x"d2c349bf",
   838 => x"a1c148c2",
   839 => x"ddff7178",
   840 => x"86c487e6",
   841 => x"48d5fac0",
   842 => x"78ced2c3",
   843 => x"fac087cc",
   844 => x"c048bfd5",
   845 => x"fac080e0",
   846 => x"d2c358d9",
   847 => x"c148bfca",
   848 => x"ced2c380",
   849 => x"0e952758",
   850 => x"97bf0000",
   851 => x"029d4dbf",
   852 => x"c387e3c2",
   853 => x"c202ade5",
   854 => x"fac087dc",
   855 => x"cb4bbfd5",
   856 => x"4c1149a3",
   857 => x"c105accf",
   858 => x"497587d2",
   859 => x"89c199df",
   860 => x"dac391cd",
   861 => x"a3c181de",
   862 => x"c351124a",
   863 => x"51124aa3",
   864 => x"124aa3c5",
   865 => x"4aa3c751",
   866 => x"a3c95112",
   867 => x"ce51124a",
   868 => x"51124aa3",
   869 => x"124aa3d0",
   870 => x"4aa3d251",
   871 => x"a3d45112",
   872 => x"d651124a",
   873 => x"51124aa3",
   874 => x"124aa3d8",
   875 => x"4aa3dc51",
   876 => x"a3de5112",
   877 => x"c151124a",
   878 => x"87fac07e",
   879 => x"99c84974",
   880 => x"87ebc005",
   881 => x"99d04974",
   882 => x"dc87d105",
   883 => x"cbc00266",
   884 => x"dc497387",
   885 => x"98700f66",
   886 => x"87d3c002",
   887 => x"c6c0056e",
   888 => x"dedac387",
   889 => x"c050c048",
   890 => x"48bfd5fa",
   891 => x"c387e1c2",
   892 => x"c048ebda",
   893 => x"dac37e50",
   894 => x"c349bfda",
   895 => x"4abfcad2",
   896 => x"fb04aa71",
   897 => x"dec387f6",
   898 => x"c005bffb",
   899 => x"dac387c8",
   900 => x"c102bfd6",
   901 => x"d2c387f8",
   902 => x"e749bfc6",
   903 => x"497087f0",
   904 => x"59cad2c3",
   905 => x"c348a6c4",
   906 => x"78bfc6d2",
   907 => x"bfd6dac3",
   908 => x"87d8c002",
   909 => x"cf4966c4",
   910 => x"f8ffffff",
   911 => x"c002a999",
   912 => x"4cc087c5",
   913 => x"c187e1c0",
   914 => x"87dcc04c",
   915 => x"cf4966c4",
   916 => x"a999f8ff",
   917 => x"87c8c002",
   918 => x"c048a6c8",
   919 => x"87c5c078",
   920 => x"c148a6c8",
   921 => x"4c66c878",
   922 => x"c0059c74",
   923 => x"66c487e0",
   924 => x"c389c249",
   925 => x"4abfceda",
   926 => x"e7dec391",
   927 => x"d2c34abf",
   928 => x"a17248c2",
   929 => x"cad2c378",
   930 => x"f978c048",
   931 => x"48c087de",
   932 => x"f1e58ef4",
   933 => x"00000087",
   934 => x"ffffff00",
   935 => x"000ea5ff",
   936 => x"000eae00",
   937 => x"54414600",
   938 => x"20203233",
   939 => x"41460020",
   940 => x"20363154",
   941 => x"1e002020",
   942 => x"bfc0dfc3",
   943 => x"05a8dd48",
   944 => x"c2c187c9",
   945 => x"497087fe",
   946 => x"ff87c84a",
   947 => x"ffc348d4",
   948 => x"724a6878",
   949 => x"1e4f2648",
   950 => x"bfc0dfc3",
   951 => x"05a8dd48",
   952 => x"c2c187c6",
   953 => x"87d987ca",
   954 => x"c348d4ff",
   955 => x"d0ff78ff",
   956 => x"78e1c848",
   957 => x"d448d4ff",
   958 => x"ffdec378",
   959 => x"bfd4ff48",
   960 => x"1e4f2650",
   961 => x"c048d0ff",
   962 => x"4f2678e0",
   963 => x"87e7fe1e",
   964 => x"02994970",
   965 => x"fbc087c6",
   966 => x"87f105a9",
   967 => x"4f264871",
   968 => x"5c5b5e0e",
   969 => x"c04b710e",
   970 => x"87cbfe4c",
   971 => x"02994970",
   972 => x"c087f9c0",
   973 => x"c002a9ec",
   974 => x"fbc087f2",
   975 => x"ebc002a9",
   976 => x"b766cc87",
   977 => x"87c703ac",
   978 => x"c20266d0",
   979 => x"71537187",
   980 => x"87c20299",
   981 => x"defd84c1",
   982 => x"99497087",
   983 => x"c087cd02",
   984 => x"c702a9ec",
   985 => x"a9fbc087",
   986 => x"87d5ff05",
   987 => x"c30266d0",
   988 => x"7b97c087",
   989 => x"05a9ecc0",
   990 => x"4a7487c4",
   991 => x"4a7487c5",
   992 => x"728a0ac0",
   993 => x"2687c248",
   994 => x"264c264d",
   995 => x"1e4f264b",
   996 => x"7087e4fc",
   997 => x"b7f0c049",
   998 => x"87ca04a9",
   999 => x"a9b7f9c0",
  1000 => x"c087c301",
  1001 => x"c1c189f0",
  1002 => x"ca04a9b7",
  1003 => x"b7dac187",
  1004 => x"87c301a9",
  1005 => x"7189f7c0",
  1006 => x"0e4f2648",
  1007 => x"0e5c5b5e",
  1008 => x"d4ff4a71",
  1009 => x"c049724c",
  1010 => x"4b7087ea",
  1011 => x"87c2029b",
  1012 => x"d0ff8bc1",
  1013 => x"78c5c848",
  1014 => x"737cd5c1",
  1015 => x"c131c649",
  1016 => x"bf97e1ec",
  1017 => x"b071484a",
  1018 => x"d0ff7c70",
  1019 => x"7378c448",
  1020 => x"87d5fe48",
  1021 => x"5c5b5e0e",
  1022 => x"86f40e5d",
  1023 => x"a6c44c71",
  1024 => x"c878c048",
  1025 => x"976e7ea4",
  1026 => x"c1c149bf",
  1027 => x"87dd05a9",
  1028 => x"9749a4c9",
  1029 => x"d2c14969",
  1030 => x"87d105a9",
  1031 => x"9749a4ca",
  1032 => x"c3c14969",
  1033 => x"87c505a9",
  1034 => x"e1c248df",
  1035 => x"87e7fa87",
  1036 => x"c3c14bc0",
  1037 => x"49bf97d3",
  1038 => x"cf04a9c0",
  1039 => x"87ccfb87",
  1040 => x"c3c183c1",
  1041 => x"49bf97d3",
  1042 => x"87f106ab",
  1043 => x"97d3c3c1",
  1044 => x"87cf02bf",
  1045 => x"7087e0f9",
  1046 => x"c6029949",
  1047 => x"a9ecc087",
  1048 => x"c087f105",
  1049 => x"87cff94b",
  1050 => x"caf94d70",
  1051 => x"58a6cc87",
  1052 => x"7087c4f9",
  1053 => x"6e83c14a",
  1054 => x"ad49bf97",
  1055 => x"c087c702",
  1056 => x"c005adff",
  1057 => x"a4c987ea",
  1058 => x"49699749",
  1059 => x"02a966c8",
  1060 => x"c04887c7",
  1061 => x"d705a8ff",
  1062 => x"49a4ca87",
  1063 => x"aa496997",
  1064 => x"c087c602",
  1065 => x"c705aaff",
  1066 => x"48a6c487",
  1067 => x"87d378c1",
  1068 => x"02adecc0",
  1069 => x"fbc087c6",
  1070 => x"87c705ad",
  1071 => x"a6c44bc0",
  1072 => x"c478c148",
  1073 => x"dcfe0266",
  1074 => x"87f7f887",
  1075 => x"8ef44873",
  1076 => x"0087f4fa",
  1077 => x"5c5b5e0e",
  1078 => x"711e0e5d",
  1079 => x"4bd4ff4d",
  1080 => x"dfc31e75",
  1081 => x"dfff49c4",
  1082 => x"86c487f7",
  1083 => x"c4029870",
  1084 => x"dfc387cb",
  1085 => x"754cbfcc",
  1086 => x"87fffa49",
  1087 => x"c005a8de",
  1088 => x"497587eb",
  1089 => x"87daf7c0",
  1090 => x"db029870",
  1091 => x"e8e3c387",
  1092 => x"e1c01ebf",
  1093 => x"e9f4c049",
  1094 => x"c186c487",
  1095 => x"c048e1ec",
  1096 => x"f4e3c350",
  1097 => x"87ecfe49",
  1098 => x"d2c348c1",
  1099 => x"48d0ff87",
  1100 => x"c178c5c8",
  1101 => x"4ac07bd6",
  1102 => x"1149a275",
  1103 => x"cb82c17b",
  1104 => x"f304aab7",
  1105 => x"c34acc87",
  1106 => x"82c17bff",
  1107 => x"aab7e0c0",
  1108 => x"ff87f404",
  1109 => x"78c448d0",
  1110 => x"c87bffc3",
  1111 => x"d3c178c5",
  1112 => x"c47bc17b",
  1113 => x"029c7478",
  1114 => x"c387c0c2",
  1115 => x"c87eced2",
  1116 => x"c08c4dc0",
  1117 => x"c603acb7",
  1118 => x"a4c0c887",
  1119 => x"c84cc04d",
  1120 => x"dc05adc0",
  1121 => x"ffdec387",
  1122 => x"d049bf97",
  1123 => x"87d10299",
  1124 => x"dfc31ec0",
  1125 => x"dde049c4",
  1126 => x"7086c487",
  1127 => x"eec04a49",
  1128 => x"ced2c387",
  1129 => x"c4dfc31e",
  1130 => x"87cae049",
  1131 => x"497086c4",
  1132 => x"48d0ff4a",
  1133 => x"c178c5c8",
  1134 => x"976e7bd4",
  1135 => x"486e7bbf",
  1136 => x"7e7080c1",
  1137 => x"ff058dc1",
  1138 => x"d0ff87f0",
  1139 => x"7278c448",
  1140 => x"87c5059a",
  1141 => x"e6c048c0",
  1142 => x"c31ec187",
  1143 => x"ff49c4df",
  1144 => x"c487f9dd",
  1145 => x"059c7486",
  1146 => x"ff87c0fe",
  1147 => x"c5c848d0",
  1148 => x"7bd3c178",
  1149 => x"78c47bc0",
  1150 => x"c2c048c1",
  1151 => x"2648c087",
  1152 => x"4c264d26",
  1153 => x"4f264b26",
  1154 => x"5c5b5e0e",
  1155 => x"711e0e5d",
  1156 => x"4d4cc04b",
  1157 => x"e8c004ab",
  1158 => x"f4ffc087",
  1159 => x"029d751e",
  1160 => x"4ac087c4",
  1161 => x"4ac187c2",
  1162 => x"d0ea4972",
  1163 => x"7086c487",
  1164 => x"6e84c17e",
  1165 => x"7387c205",
  1166 => x"7385c14c",
  1167 => x"d8ff06ac",
  1168 => x"26486e87",
  1169 => x"0e87f9fe",
  1170 => x"0e5c5b5e",
  1171 => x"66cc4b71",
  1172 => x"4c87d802",
  1173 => x"028cf0c0",
  1174 => x"4a7487d8",
  1175 => x"d1028ac1",
  1176 => x"cd028a87",
  1177 => x"c9028a87",
  1178 => x"7387d187",
  1179 => x"87e4f949",
  1180 => x"1e7487ca",
  1181 => x"ffc14973",
  1182 => x"86c487e9",
  1183 => x"0e87c3fe",
  1184 => x"5d5c5b5e",
  1185 => x"4c711e0e",
  1186 => x"c391de49",
  1187 => x"714decdf",
  1188 => x"026d9785",
  1189 => x"c387dcc1",
  1190 => x"4abfd8df",
  1191 => x"49728274",
  1192 => x"7087e5fd",
  1193 => x"c0026e7e",
  1194 => x"dfc387f2",
  1195 => x"4a6e4be0",
  1196 => x"f7fe49cb",
  1197 => x"4b7487f2",
  1198 => x"ecc193cb",
  1199 => x"83c483f1",
  1200 => x"7bf7cbc1",
  1201 => x"ccc14974",
  1202 => x"7b7587c5",
  1203 => x"97e2ecc1",
  1204 => x"c31e49bf",
  1205 => x"fd49e0df",
  1206 => x"86c487ed",
  1207 => x"cbc14974",
  1208 => x"49c087ed",
  1209 => x"87cccdc1",
  1210 => x"48c0dfc3",
  1211 => x"49c178c0",
  1212 => x"2687cfdd",
  1213 => x"4c87c9fc",
  1214 => x"6964616f",
  1215 => x"2e2e676e",
  1216 => x"5e0e002e",
  1217 => x"710e5c5b",
  1218 => x"dfc34a4b",
  1219 => x"7282bfd8",
  1220 => x"87f4fb49",
  1221 => x"029c4c70",
  1222 => x"e54987c4",
  1223 => x"dfc387e7",
  1224 => x"78c048d8",
  1225 => x"d9dc49c1",
  1226 => x"87d6fb87",
  1227 => x"5c5b5e0e",
  1228 => x"86f40e5d",
  1229 => x"4dced2c3",
  1230 => x"a6c44cc0",
  1231 => x"c378c048",
  1232 => x"49bfd8df",
  1233 => x"c106a9c0",
  1234 => x"d2c387c1",
  1235 => x"029848ce",
  1236 => x"c087f8c0",
  1237 => x"c81ef4ff",
  1238 => x"87c70266",
  1239 => x"c048a6c4",
  1240 => x"c487c578",
  1241 => x"78c148a6",
  1242 => x"e54966c4",
  1243 => x"86c487cf",
  1244 => x"84c14d70",
  1245 => x"c14866c4",
  1246 => x"58a6c880",
  1247 => x"bfd8dfc3",
  1248 => x"c603ac49",
  1249 => x"059d7587",
  1250 => x"c087c8ff",
  1251 => x"029d754c",
  1252 => x"c087e0c3",
  1253 => x"c81ef4ff",
  1254 => x"87c70266",
  1255 => x"c048a6cc",
  1256 => x"cc87c578",
  1257 => x"78c148a6",
  1258 => x"e44966cc",
  1259 => x"86c487cf",
  1260 => x"026e7e70",
  1261 => x"6e87e9c2",
  1262 => x"9781cb49",
  1263 => x"99d04969",
  1264 => x"87d6c102",
  1265 => x"4ac2ccc1",
  1266 => x"91cb4974",
  1267 => x"81f1ecc1",
  1268 => x"81c87972",
  1269 => x"7451ffc3",
  1270 => x"c391de49",
  1271 => x"714decdf",
  1272 => x"97c1c285",
  1273 => x"49a5c17d",
  1274 => x"c351e0c0",
  1275 => x"bf97deda",
  1276 => x"c187d202",
  1277 => x"4ba5c284",
  1278 => x"4adedac3",
  1279 => x"f2fe49db",
  1280 => x"dbc187e6",
  1281 => x"49a5cd87",
  1282 => x"84c151c0",
  1283 => x"6e4ba5c2",
  1284 => x"fe49cb4a",
  1285 => x"c187d1f2",
  1286 => x"c9c187c6",
  1287 => x"49744aff",
  1288 => x"ecc191cb",
  1289 => x"797281f1",
  1290 => x"97dedac3",
  1291 => x"87d802bf",
  1292 => x"91de4974",
  1293 => x"dfc384c1",
  1294 => x"83714bec",
  1295 => x"4adedac3",
  1296 => x"f1fe49dd",
  1297 => x"87d887e2",
  1298 => x"93de4b74",
  1299 => x"83ecdfc3",
  1300 => x"c049a3cb",
  1301 => x"7384c151",
  1302 => x"49cb4a6e",
  1303 => x"87c8f1fe",
  1304 => x"c14866c4",
  1305 => x"58a6c880",
  1306 => x"c003acc7",
  1307 => x"056e87c5",
  1308 => x"7487e0fc",
  1309 => x"f68ef448",
  1310 => x"731e87c6",
  1311 => x"494b711e",
  1312 => x"ecc191cb",
  1313 => x"a1c881f1",
  1314 => x"e1ecc14a",
  1315 => x"c9501248",
  1316 => x"c3c14aa1",
  1317 => x"501248d3",
  1318 => x"ecc181ca",
  1319 => x"501148e2",
  1320 => x"97e2ecc1",
  1321 => x"c01e49bf",
  1322 => x"87dbf649",
  1323 => x"48c0dfc3",
  1324 => x"49c178de",
  1325 => x"2687cbd6",
  1326 => x"1e87c9f5",
  1327 => x"cb494a71",
  1328 => x"f1ecc191",
  1329 => x"1181c881",
  1330 => x"c4dfc348",
  1331 => x"d8dfc358",
  1332 => x"c178c048",
  1333 => x"87ead549",
  1334 => x"c01e4f26",
  1335 => x"d3c5c149",
  1336 => x"1e4f2687",
  1337 => x"d2029971",
  1338 => x"c6eec187",
  1339 => x"f750c048",
  1340 => x"fbd2c180",
  1341 => x"eaecc140",
  1342 => x"c187ce78",
  1343 => x"c148c2ee",
  1344 => x"fc78e3ec",
  1345 => x"dad3c180",
  1346 => x"0e4f2678",
  1347 => x"0e5c5b5e",
  1348 => x"cb4a4c71",
  1349 => x"f1ecc192",
  1350 => x"49a2c882",
  1351 => x"974ba2c9",
  1352 => x"971e4b6b",
  1353 => x"ca1e4969",
  1354 => x"c0491282",
  1355 => x"c087f3e5",
  1356 => x"87ced449",
  1357 => x"c2c14974",
  1358 => x"8ef887d5",
  1359 => x"1e87c3f3",
  1360 => x"4b711e73",
  1361 => x"87c3ff49",
  1362 => x"fefe4973",
  1363 => x"87f4f287",
  1364 => x"711e731e",
  1365 => x"4aa3c64b",
  1366 => x"c187db02",
  1367 => x"87d6028a",
  1368 => x"dac1028a",
  1369 => x"c0028a87",
  1370 => x"028a87fc",
  1371 => x"8a87e1c0",
  1372 => x"c187cb02",
  1373 => x"49c787db",
  1374 => x"c187c0fd",
  1375 => x"dfc387de",
  1376 => x"c102bfd8",
  1377 => x"c14887cb",
  1378 => x"dcdfc388",
  1379 => x"87c1c158",
  1380 => x"bfdcdfc3",
  1381 => x"87f9c002",
  1382 => x"bfd8dfc3",
  1383 => x"c380c148",
  1384 => x"c058dcdf",
  1385 => x"dfc387eb",
  1386 => x"c649bfd8",
  1387 => x"dcdfc389",
  1388 => x"a9b7c059",
  1389 => x"c387da03",
  1390 => x"c048d8df",
  1391 => x"c387d278",
  1392 => x"02bfdcdf",
  1393 => x"dfc387cb",
  1394 => x"c648bfd8",
  1395 => x"dcdfc380",
  1396 => x"d149c058",
  1397 => x"497387ec",
  1398 => x"87f3ffc0",
  1399 => x"1e87e5f0",
  1400 => x"4b711e73",
  1401 => x"48c0dfc3",
  1402 => x"49c078dd",
  1403 => x"7387d3d1",
  1404 => x"daffc049",
  1405 => x"87ccf087",
  1406 => x"5c5b5e0e",
  1407 => x"cc4c710e",
  1408 => x"4b741e66",
  1409 => x"ecc193cb",
  1410 => x"a3c483f1",
  1411 => x"fe496a4a",
  1412 => x"c187e5ea",
  1413 => x"c87bfad1",
  1414 => x"66d449a3",
  1415 => x"49a3c951",
  1416 => x"ca5166d8",
  1417 => x"66dc49a3",
  1418 => x"d5ef2651",
  1419 => x"5b5e0e87",
  1420 => x"ff0e5d5c",
  1421 => x"a6dc86cc",
  1422 => x"48a6c859",
  1423 => x"80c478c0",
  1424 => x"7866c8c1",
  1425 => x"78c180c4",
  1426 => x"78c180c4",
  1427 => x"48dcdfc3",
  1428 => x"dfc378c1",
  1429 => x"de48bfc0",
  1430 => x"87cb05a8",
  1431 => x"7087cdf3",
  1432 => x"59a6cc49",
  1433 => x"e187d6ce",
  1434 => x"dfe287ed",
  1435 => x"87c7e187",
  1436 => x"fbc04c70",
  1437 => x"d8c102ac",
  1438 => x"0566d887",
  1439 => x"c087cac1",
  1440 => x"1ec11e1e",
  1441 => x"1ee4eec1",
  1442 => x"ebfd49c0",
  1443 => x"c086d087",
  1444 => x"d902acfb",
  1445 => x"66c4c187",
  1446 => x"6a82c44a",
  1447 => x"7481c749",
  1448 => x"d81ec151",
  1449 => x"c8496a1e",
  1450 => x"87f4e181",
  1451 => x"c8c186c8",
  1452 => x"a8c04866",
  1453 => x"c887c701",
  1454 => x"78c148a6",
  1455 => x"c8c187ce",
  1456 => x"88c14866",
  1457 => x"c358a6d0",
  1458 => x"87c0e187",
  1459 => x"c248a6d0",
  1460 => x"029c7478",
  1461 => x"c887e2cc",
  1462 => x"ccc14866",
  1463 => x"cc03a866",
  1464 => x"a6c487d7",
  1465 => x"d878c048",
  1466 => x"ff78c080",
  1467 => x"7087c8df",
  1468 => x"4866d84c",
  1469 => x"c605a8dd",
  1470 => x"48a6dc87",
  1471 => x"c17866d8",
  1472 => x"c005acd0",
  1473 => x"deff87eb",
  1474 => x"deff87ed",
  1475 => x"4c7087e9",
  1476 => x"05acecc0",
  1477 => x"dfff87c6",
  1478 => x"4c7087f2",
  1479 => x"05acd0c1",
  1480 => x"66d487c8",
  1481 => x"d880c148",
  1482 => x"d0c158a6",
  1483 => x"d5ff02ac",
  1484 => x"a6e0c087",
  1485 => x"7866d848",
  1486 => x"c04866dc",
  1487 => x"05a866e0",
  1488 => x"c087c8ca",
  1489 => x"c048a6e4",
  1490 => x"c080c478",
  1491 => x"c04d7478",
  1492 => x"c9028dfb",
  1493 => x"8dc987ce",
  1494 => x"c287db02",
  1495 => x"f7c1028d",
  1496 => x"028dc987",
  1497 => x"c487d1c4",
  1498 => x"c2c1028d",
  1499 => x"028dc187",
  1500 => x"c887c5c4",
  1501 => x"66c887e8",
  1502 => x"c191cb49",
  1503 => x"c48166c4",
  1504 => x"7e6a4aa1",
  1505 => x"e8c11e71",
  1506 => x"66c448f5",
  1507 => x"4aa1cc49",
  1508 => x"aa714120",
  1509 => x"87f8ff05",
  1510 => x"49265110",
  1511 => x"79dfd7c1",
  1512 => x"87e8ddff",
  1513 => x"e8c04c70",
  1514 => x"78c148a6",
  1515 => x"c487f5c7",
  1516 => x"f0c048a6",
  1517 => x"fedbff78",
  1518 => x"c04c7087",
  1519 => x"c002acec",
  1520 => x"a6c887c3",
  1521 => x"acecc05c",
  1522 => x"ff87cd02",
  1523 => x"7087e8db",
  1524 => x"acecc04c",
  1525 => x"87f3ff05",
  1526 => x"02acecc0",
  1527 => x"ff87c4c0",
  1528 => x"c487d4db",
  1529 => x"66d81e66",
  1530 => x"66d81e49",
  1531 => x"eec11e49",
  1532 => x"66d81ee4",
  1533 => x"87c0f849",
  1534 => x"1eca1ec0",
  1535 => x"4966e0c0",
  1536 => x"dcc191cb",
  1537 => x"a6d88166",
  1538 => x"78a1c448",
  1539 => x"49bf66d8",
  1540 => x"87ccdcff",
  1541 => x"b7c086d8",
  1542 => x"cbc106a8",
  1543 => x"de1ec187",
  1544 => x"bf66c81e",
  1545 => x"f7dbff49",
  1546 => x"7086c887",
  1547 => x"08c04849",
  1548 => x"a6ecc088",
  1549 => x"a8b7c058",
  1550 => x"87ecc006",
  1551 => x"4866e8c0",
  1552 => x"03a8b7dd",
  1553 => x"6e87e1c0",
  1554 => x"e8c049bf",
  1555 => x"e0c08166",
  1556 => x"66e8c051",
  1557 => x"6e81c149",
  1558 => x"c1c281bf",
  1559 => x"66e8c051",
  1560 => x"6e81c249",
  1561 => x"51c081bf",
  1562 => x"c14866d0",
  1563 => x"58a6d480",
  1564 => x"c180d848",
  1565 => x"87ecc478",
  1566 => x"87d3dcff",
  1567 => x"58a6ecc0",
  1568 => x"87cbdcff",
  1569 => x"58a6f0c0",
  1570 => x"05a8ecc0",
  1571 => x"a687c9c0",
  1572 => x"66e8c048",
  1573 => x"87c4c078",
  1574 => x"87dbd8ff",
  1575 => x"cb4966c8",
  1576 => x"66c4c191",
  1577 => x"c8807148",
  1578 => x"66c458a6",
  1579 => x"c482c84a",
  1580 => x"81ca4966",
  1581 => x"5166e8c0",
  1582 => x"4966ecc0",
  1583 => x"e8c081c1",
  1584 => x"48c18966",
  1585 => x"49703071",
  1586 => x"977189c1",
  1587 => x"c8e3c37a",
  1588 => x"e8c049bf",
  1589 => x"6a972966",
  1590 => x"9871484a",
  1591 => x"58a6f4c0",
  1592 => x"c44966c4",
  1593 => x"c07e6981",
  1594 => x"dc4866e0",
  1595 => x"c002a866",
  1596 => x"a6dc87c8",
  1597 => x"c078c048",
  1598 => x"a6dc87c5",
  1599 => x"dc78c148",
  1600 => x"e0c01e66",
  1601 => x"4966c81e",
  1602 => x"87d4d8ff",
  1603 => x"4c7086c8",
  1604 => x"06acb7c0",
  1605 => x"6e87d6c1",
  1606 => x"70807448",
  1607 => x"49e0c07e",
  1608 => x"4b6e8974",
  1609 => x"4af2e8c1",
  1610 => x"fbddfe71",
  1611 => x"c2486e87",
  1612 => x"c07e7080",
  1613 => x"c14866e4",
  1614 => x"a6e8c080",
  1615 => x"66f0c058",
  1616 => x"7081c149",
  1617 => x"c5c002a9",
  1618 => x"c04dc087",
  1619 => x"4dc187c2",
  1620 => x"a4c21e75",
  1621 => x"48e0c049",
  1622 => x"49708871",
  1623 => x"4966c81e",
  1624 => x"87fcd6ff",
  1625 => x"b7c086c8",
  1626 => x"c6ff01a8",
  1627 => x"66e4c087",
  1628 => x"87d3c002",
  1629 => x"c94966c4",
  1630 => x"66e4c081",
  1631 => x"4866c451",
  1632 => x"78cbd4c1",
  1633 => x"c487cec0",
  1634 => x"81c94966",
  1635 => x"66c451c2",
  1636 => x"ffd4c148",
  1637 => x"a6e8c078",
  1638 => x"c078c148",
  1639 => x"d5ff87c6",
  1640 => x"4c7087ea",
  1641 => x"0266e8c0",
  1642 => x"c887f5c0",
  1643 => x"66cc4866",
  1644 => x"cbc004a8",
  1645 => x"4866c887",
  1646 => x"a6cc80c1",
  1647 => x"87e0c058",
  1648 => x"c14866cc",
  1649 => x"58a6d088",
  1650 => x"c187d5c0",
  1651 => x"c005acc6",
  1652 => x"66d087c8",
  1653 => x"d480c148",
  1654 => x"d4ff58a6",
  1655 => x"4c7087ee",
  1656 => x"c14866d4",
  1657 => x"58a6d880",
  1658 => x"c0029c74",
  1659 => x"66c887cb",
  1660 => x"66ccc148",
  1661 => x"e9f304a8",
  1662 => x"c6d4ff87",
  1663 => x"4866c887",
  1664 => x"c003a8c7",
  1665 => x"dfc387e5",
  1666 => x"78c048dc",
  1667 => x"cb4966c8",
  1668 => x"66c4c191",
  1669 => x"4aa1c481",
  1670 => x"52c04a6a",
  1671 => x"4866c879",
  1672 => x"a6cc80c1",
  1673 => x"04a8c758",
  1674 => x"ff87dbff",
  1675 => x"dfff8ecc",
  1676 => x"203a87ce",
  1677 => x"50494400",
  1678 => x"69775320",
  1679 => x"65686374",
  1680 => x"731e0073",
  1681 => x"9b4b711e",
  1682 => x"c387c602",
  1683 => x"c048d8df",
  1684 => x"c31ec778",
  1685 => x"49bfd8df",
  1686 => x"f1ecc11e",
  1687 => x"c0dfc31e",
  1688 => x"c8ef49bf",
  1689 => x"c386cc87",
  1690 => x"49bfc0df",
  1691 => x"7387f4e9",
  1692 => x"87c8029b",
  1693 => x"49f1ecc1",
  1694 => x"87e5eec0",
  1695 => x"87c4deff",
  1696 => x"e1ecc11e",
  1697 => x"c150c048",
  1698 => x"49bfd4ee",
  1699 => x"87c4d9ff",
  1700 => x"4f2648c0",
  1701 => x"87ebc71e",
  1702 => x"e5fe49c1",
  1703 => x"eee2fe87",
  1704 => x"02987087",
  1705 => x"ebfe87cd",
  1706 => x"987087e9",
  1707 => x"c187c402",
  1708 => x"c087c24a",
  1709 => x"059a724a",
  1710 => x"1ec087ce",
  1711 => x"49e8ebc1",
  1712 => x"87fef9c0",
  1713 => x"87fe86c4",
  1714 => x"87f0e5c1",
  1715 => x"ebc11ec0",
  1716 => x"f9c049f3",
  1717 => x"1ec087ec",
  1718 => x"7087e5fe",
  1719 => x"e1f9c049",
  1720 => x"87dec387",
  1721 => x"4f268ef8",
  1722 => x"66204453",
  1723 => x"656c6961",
  1724 => x"42002e64",
  1725 => x"69746f6f",
  1726 => x"2e2e676e",
  1727 => x"c01e002e",
  1728 => x"c187fff0",
  1729 => x"f687c6de",
  1730 => x"1e4f2687",
  1731 => x"48d8dfc3",
  1732 => x"dfc378c0",
  1733 => x"78c048c0",
  1734 => x"e187f9fd",
  1735 => x"2648c087",
  1736 => x"8000004f",
  1737 => x"69784520",
  1738 => x"20800074",
  1739 => x"6b636142",
  1740 => x"0014bb00",
  1741 => x"0037ec00",
  1742 => x"00000000",
  1743 => x"000014bb",
  1744 => x"0000380a",
  1745 => x"bb000000",
  1746 => x"28000014",
  1747 => x"00000038",
  1748 => x"14bb0000",
  1749 => x"38460000",
  1750 => x"00000000",
  1751 => x"0014bb00",
  1752 => x"00386400",
  1753 => x"00000000",
  1754 => x"000014bb",
  1755 => x"00003882",
  1756 => x"bb000000",
  1757 => x"a0000014",
  1758 => x"00000038",
  1759 => x"14bb0000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00155000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00001b98",
  1766 => x"544f4f42",
  1767 => x"20202020",
  1768 => x"004d4f52",
  1769 => x"64616f4c",
  1770 => x"002e2a20",
  1771 => x"48f0fe1e",
  1772 => x"09cd78c0",
  1773 => x"4f260979",
  1774 => x"f0fe1e1e",
  1775 => x"26487ebf",
  1776 => x"fe1e4f26",
  1777 => x"78c148f0",
  1778 => x"fe1e4f26",
  1779 => x"78c048f0",
  1780 => x"711e4f26",
  1781 => x"5252c04a",
  1782 => x"5e0e4f26",
  1783 => x"0e5d5c5b",
  1784 => x"4d7186f4",
  1785 => x"c17e6d97",
  1786 => x"6c974ca5",
  1787 => x"58a6c848",
  1788 => x"66c4486e",
  1789 => x"87c505a8",
  1790 => x"e6c048ff",
  1791 => x"87caff87",
  1792 => x"9749a5c2",
  1793 => x"a3714b6c",
  1794 => x"4b6b974b",
  1795 => x"6e7e6c97",
  1796 => x"c880c148",
  1797 => x"98c758a6",
  1798 => x"7058a6cc",
  1799 => x"e1fe7c97",
  1800 => x"f4487387",
  1801 => x"264d268e",
  1802 => x"264b264c",
  1803 => x"5b5e0e4f",
  1804 => x"86f40e5c",
  1805 => x"66d84c71",
  1806 => x"9affc34a",
  1807 => x"974ba4c2",
  1808 => x"a173496c",
  1809 => x"97517249",
  1810 => x"486e7e6c",
  1811 => x"a6c880c1",
  1812 => x"cc98c758",
  1813 => x"547058a6",
  1814 => x"caff8ef4",
  1815 => x"fd1e1e87",
  1816 => x"bfe087e8",
  1817 => x"e0c0494a",
  1818 => x"cb0299c0",
  1819 => x"c31e7287",
  1820 => x"fe49fee2",
  1821 => x"86c487f7",
  1822 => x"7087fdfc",
  1823 => x"87c2fd7e",
  1824 => x"1e4f2626",
  1825 => x"49fee2c3",
  1826 => x"c187c7fd",
  1827 => x"fc49ddf1",
  1828 => x"c8c487da",
  1829 => x"1e4f2687",
  1830 => x"c848d0ff",
  1831 => x"d4ff78e1",
  1832 => x"c478c548",
  1833 => x"87c30266",
  1834 => x"c878e0c3",
  1835 => x"87c60266",
  1836 => x"c348d4ff",
  1837 => x"d4ff78f0",
  1838 => x"ff787148",
  1839 => x"e1c848d0",
  1840 => x"78e0c078",
  1841 => x"5e0e4f26",
  1842 => x"710e5c5b",
  1843 => x"fee2c34c",
  1844 => x"87c6fc49",
  1845 => x"b7c04a70",
  1846 => x"e3c204aa",
  1847 => x"aae0c387",
  1848 => x"c187c905",
  1849 => x"c148d0f6",
  1850 => x"87d4c278",
  1851 => x"05aaf0c3",
  1852 => x"f6c187c9",
  1853 => x"78c148cc",
  1854 => x"c187f5c1",
  1855 => x"02bfd0f6",
  1856 => x"4b7287c7",
  1857 => x"c2b3c0c2",
  1858 => x"744b7287",
  1859 => x"87d1059c",
  1860 => x"bfccf6c1",
  1861 => x"d0f6c11e",
  1862 => x"49721ebf",
  1863 => x"c887f8fd",
  1864 => x"ccf6c186",
  1865 => x"e0c002bf",
  1866 => x"c4497387",
  1867 => x"c19129b7",
  1868 => x"7381ecf7",
  1869 => x"c29acf4a",
  1870 => x"7248c192",
  1871 => x"ff4a7030",
  1872 => x"694872ba",
  1873 => x"db797098",
  1874 => x"c4497387",
  1875 => x"c19129b7",
  1876 => x"7381ecf7",
  1877 => x"c29acf4a",
  1878 => x"7248c392",
  1879 => x"484a7030",
  1880 => x"7970b069",
  1881 => x"48d0f6c1",
  1882 => x"f6c178c0",
  1883 => x"78c048cc",
  1884 => x"49fee2c3",
  1885 => x"7087e3f9",
  1886 => x"aab7c04a",
  1887 => x"87ddfd03",
  1888 => x"87c248c0",
  1889 => x"4c264d26",
  1890 => x"4f264b26",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"494a711e",
  1894 => x"2687ebfc",
  1895 => x"4ac01e4f",
  1896 => x"91c44972",
  1897 => x"81ecf7c1",
  1898 => x"82c179c0",
  1899 => x"04aab7d0",
  1900 => x"4f2687ee",
  1901 => x"5c5b5e0e",
  1902 => x"4d710e5d",
  1903 => x"7587cbf8",
  1904 => x"2ab7c44a",
  1905 => x"ecf7c192",
  1906 => x"cf4c7582",
  1907 => x"6a94c29c",
  1908 => x"2b744b49",
  1909 => x"48c29bc3",
  1910 => x"4c703074",
  1911 => x"4874bcff",
  1912 => x"7a709871",
  1913 => x"7387dbf7",
  1914 => x"87d8fe48",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"00000000",
  1927 => x"00000000",
  1928 => x"00000000",
  1929 => x"00000000",
  1930 => x"00000000",
  1931 => x"48d0ff1e",
  1932 => x"7178e1c8",
  1933 => x"08d4ff48",
  1934 => x"4866c478",
  1935 => x"7808d4ff",
  1936 => x"711e4f26",
  1937 => x"4966c44a",
  1938 => x"ff49721e",
  1939 => x"d0ff87de",
  1940 => x"78e0c048",
  1941 => x"1e4f2626",
  1942 => x"4b711e73",
  1943 => x"1e4966c8",
  1944 => x"e0c14a73",
  1945 => x"d9ff49a2",
  1946 => x"87c42687",
  1947 => x"4c264d26",
  1948 => x"4f264b26",
  1949 => x"4ad4ff1e",
  1950 => x"ff7affc3",
  1951 => x"e1c848d0",
  1952 => x"c37ade78",
  1953 => x"7abfc8e3",
  1954 => x"28c84849",
  1955 => x"48717a70",
  1956 => x"7a7028d0",
  1957 => x"28d84871",
  1958 => x"d0ff7a70",
  1959 => x"78e0c048",
  1960 => x"5e0e4f26",
  1961 => x"0e5d5c5b",
  1962 => x"e3c34c71",
  1963 => x"4b4dbfc8",
  1964 => x"66d02b74",
  1965 => x"d483c19b",
  1966 => x"c204ab66",
  1967 => x"744bc087",
  1968 => x"4966d04a",
  1969 => x"b9ff3172",
  1970 => x"48739975",
  1971 => x"4a703072",
  1972 => x"c3b07148",
  1973 => x"fe58cce3",
  1974 => x"4d2687da",
  1975 => x"4b264c26",
  1976 => x"5e0e4f26",
  1977 => x"0e5d5c5b",
  1978 => x"c34c711e",
  1979 => x"c04bcce3",
  1980 => x"49f4c04a",
  1981 => x"87cdc7fe",
  1982 => x"e3c31e74",
  1983 => x"e7fe49cc",
  1984 => x"86c487df",
  1985 => x"02994970",
  1986 => x"c487eac0",
  1987 => x"1e4da61e",
  1988 => x"49cce3c3",
  1989 => x"87e3eefe",
  1990 => x"987086c8",
  1991 => x"7587d602",
  1992 => x"ebfdc14a",
  1993 => x"fe4bc449",
  1994 => x"7087ffc4",
  1995 => x"87ca0298",
  1996 => x"edc048c0",
  1997 => x"c048c087",
  1998 => x"f3c087e8",
  1999 => x"87c4c187",
  2000 => x"c8029870",
  2001 => x"87fcc087",
  2002 => x"f8059870",
  2003 => x"ece3c387",
  2004 => x"87cc02bf",
  2005 => x"48c8e3c3",
  2006 => x"bfece3c3",
  2007 => x"87d4fc78",
  2008 => x"262648c1",
  2009 => x"264c264d",
  2010 => x"5b4f264b",
  2011 => x"00435241",
  2012 => x"c31ec01e",
  2013 => x"fe49cce3",
  2014 => x"c387d9eb",
  2015 => x"c048e4e3",
  2016 => x"4f262678",
  2017 => x"5c5b5e0e",
  2018 => x"86f40e5d",
  2019 => x"c048a6c4",
  2020 => x"e4e3c378",
  2021 => x"b7c348bf",
  2022 => x"87d103a8",
  2023 => x"bfe4e3c3",
  2024 => x"c380c148",
  2025 => x"c058e8e3",
  2026 => x"e2c648fb",
  2027 => x"cce3c387",
  2028 => x"daf0fe49",
  2029 => x"c34c7087",
  2030 => x"4abfe4e3",
  2031 => x"d8028ac3",
  2032 => x"028ac187",
  2033 => x"8a87cbc5",
  2034 => x"87f6c202",
  2035 => x"cdc1028a",
  2036 => x"c3028a87",
  2037 => x"e1c587e2",
  2038 => x"754dc087",
  2039 => x"c292c44a",
  2040 => x"c382edc5",
  2041 => x"7548e0e3",
  2042 => x"6e7e7080",
  2043 => x"494bbf97",
  2044 => x"c1486e4b",
  2045 => x"816a50a3",
  2046 => x"a6cc4811",
  2047 => x"02ac7058",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
